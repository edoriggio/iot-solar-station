PK   ��Wx�D��,  ��    cirkitFile.json�]o�F����B}+
I2�<w��1��mL/z/|
d�l#Kg�:��1��7���*UɊ7$�g�@۪�
>|��Hf�zl���/����o�������'*��~j�_����뫯�����⯏�ן�>�*g�|���o�����sח�����uYQuV��ϖ��}��K_��pW�~�r}�R[pR3h-��W3h-�E�f�Zp�B͠����Ak�-��Ak�-��Ak�-*5�Xx��������jQ�E����������Z�Y�jOl�q]��t}�m[�e�Y����5u�Y�w˾�]��<��~��]6��Ɋ�鳺(�k]Q���+('��uJ�̖u��\�<k=U�gY��P�q)!��o�!,]`R_-���<�o߸����������\�F쉓N;W�=q��Ğ`N�Tb�Zleϧ�~�&���{`�w�jL���&�B��M0��#V�`
}W�6���Xm�)�ݱ�Sh�M��];�&�B;�&����c���N�	���N�	���N�	���N�	���N�	���N�	���N�	����Sm�)��Sm�)��Sm�) �?�ؙ�c��S�c��S�c��S�c��S�c��S�c�ڄ[�ة6��ة6��ة6��ة6���s}�,��Sm�)��Sm�)��Sm�)��Sm�)��Sm�-J}�T�`
}�T�`
}�T�`
}�T�`
}�T�`
��G}�,��Sm�)��Sm�)��Sm�)��Sm�-�>v�M0�>v�M0�>v�L|}����ۻ�3��w�����㧉'�IOO��H���jHHEBi�$=��8�iM�Hr�աcM`�6'��iDw�x����$��y���+�#,�[�X�r�vP:��q��ծ�j�#,��X�J�v#�S�-i��n�@����t��	⊍Nfn�sKZ.�,F�SN,�t�,���I�X��b�F����-j�v5V;(a�dy*8s�dʄ�G`>YX���A��'K����R��YSj���:VNy�9"��D,��dy8X?p���#0�,l�N�|�%�`������|�� �4� 0��dX?pF��#0�l� �Ί�|擭'����G`>�4��a��'�}���P��P�Qyp�������|��
�8����O6����X>�ɶ6�~���G`>ِ��`��'[	����,��d$X?p���#0�l����X>���S�~���G`>�2��`��'�}���ɡWɁ������G`>�`��`��'[�����,��dS;X?p���#0�l���?�|�B`������|R�_�?�|��`������|Rv�8����O
f���X>�I��~�:�:��� �8����Oʫ���X>�Ia�~���G`>)i��`��'�x����,����V��`��'�����,���tX?p���#0����?�|�rY`������|R���X 8���I�2�~���G`>)���`��'e�����,����X?p���#0����������|RD�8����O����X>:�7�~�n����LA�U$��K
�\IrԿ+H��K�6�88�.o_<}����k�R�!�(�d�_�i�������"_�(R�A�Pm�A�A�������0*>���P��g�h+�j�5
y�C,\��>�xTWo�K͑Is�9��9N�|�&o�n�ڬp}�Q�j3b݆6~�ujO�+9��*�'_�rd���&놈B�z���C_fU��Y(�~�j��.S�4��:�DU�'�#O�sb8P�k�\L��Tq�>$�Tyr0��G�GN|�͈!��6#��
�ʒr)#�$�|���s<򭩍YQ�8TY�nh����A5��Sc��#O��Ī�0���̉��(^?�/����đ�ޒ`u�'��O|S���2��7U�H��������� �8$��#�o�c/V������է_5��J\��������  C�.C2��71D C��C2��W1D C��C2�d� C2�d.C2�d�C�6���tD���ʢ�հ	�(Kn=Yb��m�n�%)c��n�o�%)Zc��o�p�%)�c��p�q�%)c��q��(KR�Ƅ��8�aqeI
U`q���8ʒT�1�⸇�q�%)�c��q��(KR�����x��(KRHƄ�I�M���x��(KRD���9,��,I�',��8��$E�`L�8^��8ʒρ1��x��(KR�Ƅ��M���x��(KR����,��,I!
,��8��$`�~`q���q�%��c����Q�d:�	�t�x�KXGY���0&X/aqeI6�`q<��8ʒl�1��x���)K��^l���V�;-��@U�/���n��j5�;^��Z�;�VG�A��Y��	��z�3��+����q�"�U���d��y���Ǖ�0
X��	�;�?��
�ů����j ���q�#��cV�U`�u\	s��+"a�YcV���Y
�H�[��+����q�$�U���d�*k�m�q�,hɆV�6�hk�uYВ��Ѷ�v�� z0Z�����6��d_&�dC+k�m����LhɆV���hk���В��a���&3�%Zًa��E�C6�dC+{Jl����LhɆV���hk���В���y�`���В��U���&/3�%Z�se���1�Gb6�ļM^�m�2Z���=p6���e&�dC+{�l����LhɆV�$�hk���В�쭴��&/3�%Z�#j��M^fBK6����F[��̄�lheϮ��$��̄�lheﱍ�6y�	-���jmm�2Z�����6��V4Z�h���6yYn���В��ͷ��&/3�%Z�1`��M^fBK6�R+�F[��̄�lh�惍�6y�	-��J�
mm�2Z���&�6y�	-��J-mm�2Z����(6���e&�dC+�]l����LhɆVj��hk���h+�M^V��e�M^fBK6�R3�F[��̄�lh�����6y�	-��J'mm�2Z���ZT6���e&�dC+5�L�-m�2Z����`6���e&�dC+5�l����LhɆVj��hk���В�Ԝ���&/3�%Z��g��Q���̄Vj �hk���В��2���&/3�%Z��h��M^fBK6�R[�F[��̄�lh�F����&/3�%Z��i��M^fBK6�R��F[��̄��h�_]�E����.�!+b��y���q]�y��L+be]�{\�d��u���\gZ�V�=~�볕���2_��	��x���1+��n�����Yu���9]���s�$Y����brw��^o~�x���t�����a(��ʺB�������DM��V�UЇv�QXY�-%�D��^�60y�W3��������t>E[q��}ֆ<φ!�l{�6¨��9�I���yo��M�f�ҵY���#L�f.ĺm�ҟ?�$+t�c���sޛ�uJ�̖u�=w��T�eY7CYƥۜ�kq*���)��ٞ:�J�Q��
+o��i�<ח�sܯ��Ƭ�����*�|�M�qoן��$+tN�nKǦ2��"+:�c��qQ5y?��yI�r�_�����$+gGv�n�(Ĭ���ơ/��n�,�u�t5�ʄk�d�^����f���ӪY�W�~}6;��
�w�[=6w/��Wdh3 D C��!��2��&.B�@�61B2�֣SȐ[�t!D Cn=j����B2�6�yL��Em\؆�m�n�%�,c��n�o�%�d
c��o�p�%��	c��p�q�%��c��q��(KRƄ��8�aqeI*���`q���8ʒT�1�⸇�q�%�Pc��q��(KR	����x��(KR�Ƅ�I�M���x��(KR)���9,��,Ie,��8��$� `L�8^��8ʒT�1��x��(K��Ƅ��M���x��(K�#���,��,�X,��8��$;.a�~`q���q�%��c����Q�dG�	�t�x�KXGY��?0&X/aqeIv���`q<��8ʒ�l�1��x���)K�w)�v���n6 ��	+����h�*PWV2au����U���d����h�@]-XɄ��.]G� 
X��	+��Lt"�(`�J&�<F1�uT� ��+���Ũ�*PWV2au�Q��U���d����h�@]-XɄU��$6�	-����fm��.���&�"�ċl2/Z�����6��d_&�dC+k�m����LhɆV���hk���В��a���&3�%Zًa��M6fBK6����F[��̄�lheo���6Y�	-����6y�	-���^%mm�2Z���=W6�=3z$f��y�����e&�dC+{�l����LhɆV���hk���В��I���&/3�%Z�[i��M^fBK6��G�F[��̄�lhe����6y�	-��ʞ]��I6y�	-����cmm�2Z���=�6���e&�dC+{�m�5Z�h�\�&/�m��&/3�%Zٛo��M^fBK6�Rc�F[��̄�lh�V���6y�	-��J�mm�2Z����6���e&�dC+58L�-l�2Z���Z"6���e&�dC+5Ql����LhɆVj��hk���В�Ԩ���h'��V2������
��̄�lh�f���6y�	-��J�#mm�2Z���N6���e&�dC+��l����LhɆVjj�h[��e&�dC+��l����LhɆVj��hk���В��j���&/3�%Z�9g��M^fBK6�R;�F[�*Fe>l��&/+m�2Z���Z�6���e&�dC+5m����LhɆVjK�hk���В���4�6��e&�dC+�>m����LhɆVj��hk����R�׿�E����.�!+b��y���q];��V&��δ2Q�{�����3�LT�}�Ҷu_�ː5!��c��1f���-�>v<�8�n���k�d��5���a�eCh���>���2_����ۼ:�K����$Y9�K��.g}7��D���V&j�ϴ2Q}�����3�LT��u �=뽾��t>E[q��}ֆ<φ!�l{cB�I��a9��y��Y�tmV���S���nC��	=R���g�d���y݅�-�e]p�]�<k=U�gY��P�q�ΟQ���g�dsFg�]����.���h|�q�VS������]74yǽ]�%Y9{��!,��|�,���<���51P��C�0&K��a9�/IV��K�"
1��q�ˬ��:e�/]�ò2�%Yy��o���_-�w�����W�|}}���c���z�,�nq{�xx��ǫO?��f��<����$���(�Ӑ/I�ƢV�t�A���/��O�Ki�ڣ�{�R�w�Sw�w��^��tOLm�<1�T��;�N����(��_�p��LTݜ��Sw�*��OI��� �WN0�2p�;��$��&��]{������o����R����S;��ccZ6�d��8����l�N��no9i1zߔM(r}�Ta=�[F�5�Hչ2��s�J*ۼ�'N=@��'�`ү�� m$�$G���+5A���OER%i��$ZMF̗�l��Dv�(��8[#;.X��+���7&��o<k�h4(U�5���\��yb�?�J}8K\:�Y�9��:GՑ5׹�(j�kG��b$�D�9��,ޖ�pEՃI}�[��=�O\��"ym��˼|����}VU��>Ħ�9.�S� q1�đ�h i�<yu���ڴ��z�k�I`�1q͕MdL\�5q�h�A<J\���(qu�f����)qqڗ/��g����EsߝZ��#C~�i_F^���/O�3 V��!�u��P��W�����P���+�|$�B�p��+���=�;����n��l�R��uZ��_Н���w�Q���C��!m���}p��E�z��'�>�r�c�yg������v��?�?��'G?yi�w��R!��
B!�v�H��������:h~/#�2"R�1���ڹ�w�O���!�;S8�Dd����� �n�h�'�� �[>H
c{�Q������3"� o��Rw	Y�0�nz�¼Ǟ���]hθ�{�e��w*��%�3�V����3����&���M��K�nZ�w��X
�_k�F[�̒��5�Ə�1>���r?���
���73��-�>�z���G0��@��r����(w��PnϜvҷآ��p�MN_���3����
@�:��N�W�ٿ���ͥ���a=�r���~����fD(13��[�-uH�q��������М	��!\���@���+}fb�V"�Yy�m�z �n���m��E~�[�đ�5ﻻ�`��+�~�" �}vj-�W/�{���+觞� �:�p�N����a�jV�է��ð��X=,��vW�~�8��yg�{h�6�y��Bmb�-%����\J
�����j�7�))�&��}�J
�	�~ߢ�Bm­�ר���\U�-�j|�ڢ6�B�ކۼ�R����z�Rz@�%@���`@���`@���`@���`@���`u,$����s ��s ���x��To�9 �To�9 �To�9 �To�9 �To�9 �To�9 �To��L@<��`@<��`@<��`�  ��x����x����x����x����x����x��� ��m0 ��m0 ��m0 ��m0bJO@<��`@<��`@<��`@<��`@<��p�O�6�O�6�O�6�O�6�O�6��
OK@<��`@<��`@<��`@<��p� ��z���z���c�A�'���Z�I#��E��rk�z�, E���kIǸ*{��ǧOf���ujx���.���|n������a��玷 �A������qBڃ�7�;�ڔ��;*�;�U�`uG�8{'"���#�Y�\��cTad�����nV�;+�oT-H}�5X�����|��=Reڡ:��Є�P����&�@�<�Ϩr0B�+�b�ey.Zat�&$4�,-Fk�N}���&�e�h����Є���!:��P���5���&$4�,�Gk��_���&�m h�9��Є��=#��b���&��h�Y��Є�u�!������G�)���		M([v���0!�	e�ZCt�&$4�l�Bk��S���&�m^h�y
��Є�E�!:O�P�ס5D�)`BB��@��t�&$4�lkDk��S���&�-�h�y
��Є���!||:O��yJ��S���&�m�h�y
��Є��!:O�P�O�5D�)`BB��o���<LHhBٶ�����		M([���<LHhB)�����		M(����0!�	�LZCt�&$4���@k�����S
t�R��0!�	��ZCt�&$4��%Ak��S���&��*h�y
��ЄR�!:O�PJـ5,�y
��ЄR��!:O�PJ�5D�)`BBJ�#���<LHhB)݄����		M(e��·��0���Bk��S���&�r_h�y
��ЄR��!:O�Pʬ�5D�)`BBJ�8�����		M(�����0!�	�4ZCt�&�s��/���������Ր��YC�<�U퉭7�kׯd|��Ls~ln��I�򱹉wv&�+��&��d�����ڶ��|�&6�}̚:Ƭ�޻e�ǎG
'.E�0w��+̝���%�;qe'�Kz��	�&^��^��M2wB;�ɞ�n�m�I��w��ki�̕cs�l��067��I��؜�ʎ�PI�+;~=%M������jΖ��������t>E[q �}ֆ<φ!�l{㩈7um�̍�</������/��v��ͺ�k���G���\�u�0��?u��6�܉���$s'Nv�S��"k̥��I�N��Ġ'��8�D<N2w"O�eI�N��x�\�18�wMm̊zh�\���w���w��)7��K2w'�Kz�|��%�K��$sc��%��������=���'��߮����v�fz��$��Or_}��J.��r1����Uʘs�c����{�n�,�[��Nr�㮻Z3�t2���G)�z���80}l �V}6�?H�ϓz��΋#��|۸�}�/Y�lftS�O��z�k�5}�&��dP��D��Ӂ���|Ռ����i�T/=Ur��*ϥ�fd����Lth�;&qp0��O8G���9�9�-5p�"������8.��=66��(�|7IyN�z.q:H��U8�r��e������kf��0S�`��f�m3�gf43vc�|��K������a
��2U'`�b|✒f�q3u�'�h�<�0SA1q^A3�3���>�t�ۙMQ�zk���P#8?�gLTp�1~*b'ο��N+7�S��5SAc����$B3��b`��}��k��N�e�����!���W����_��Wn�U��*�_��W���r�U�~�_��Wa�U���Um��F_��h|b��c��ΌƧF;Ah��ԧ�����ƚ����9�ΜƧN;�h��t���~����w���.~�Ǻ��.�9���n�"���w�O+����C�~�����̫���*�/��V�Ϸ9���}�_ͪ�����Ǉ���궗)\>q����ۇ{n�U���ˢ�����5�q�2����D6,����<tu�<�GJ*3�8䖱��9T������Ӫ�_n~�4g|}��x����{��?\�>.����0m�o�k&�r���Ţ(��'E�Ob���d���)P�.'�bn�P�!_�ܮ.���Uq�F�m��뢮o*V?��F��˗5�ܮ�����>��|ڠ��xv���Ub^]�uqS����9�K��bY�mWey,zV�)��[Y��P45��X����cտ}kNT��9��MA��}Y;������낶���/ٽ�|����B�=�Y���uV��O;���z��ӻ�C�&PV�X4�}�����=V2��C����|�Y�o���eY�U��˛���"ߵ�7�ے���o"nK����뛜��P�O�75��U~S�%7�}�������b�zuص�|����͔�^eȣ�5��-Å�1rr<r-w�P�w��%z�2�~\훐gS܄ʛ������n�˛���$V�U/%���X�m�^��(ϋ݉]�eW?���q˧���L��7?������ߚ�o�׿��;��:H���������O������OCs���O��_n�nۻ~��c����>��u+����?7�߆f����?����3˟�6�����{ �q���AE����;���o���=�8�:��}�����'vY��}�Cp�rM5�ׂ�xI��f�x��)v��xYD�oߘ��r�	���F�������;�b��ߔ��7с���!.p���N�C����r��˳tU��v�Z��gE�S֖<��ˮ�z��<�:�.���t��A.����@�*�?��ݕy����&U2X�3�oBQq��=�u'F���2F��w��h{�ܷ�M^{��j�*�W���G�%'��[�7��<�\Vgs��� ��;���b�����T�l3Δy���5-�.t���$=�O���|��.ۿ�E[�Όۋr�T��bߟ?�b�۹�)+��ɪ%QF����*��$�@���
�.�e��ᘕ�#P��G����>婟���T�×�-*�>���T��wyB(o"��4�~Qn7�pہ����Q�~�����o��Uκ�r�c�X�e�B�]%_�nY��|�%i|�oʗ��{�����c�ס���y|y��M���X�o�ݺ^=p�uţ��׶^Ϧ�]�?#!�=G���n��؈���O��_��<v2L2s��я�qxY(�,�������j�������_�!�$���3_ệ��W�>_�A�Y�����g������_i�Ƭ����	ksW��M=6���,]������dʅ��W�ׇ����꧵�_?�|%�+~�/��=ɧ�~���x���=�{����T3�O6;�*Hn��N(�;����7���,i˛,��R�e��Y8�?yyyXpQ��Y�����k�>���-i���"�_f�j��H
.��9G͞gvN7�p^����|��@�zA<������ �z5�3���>���-f���<�_f�j�%��=�*^Ќ���(^�n�+���w�U����=����uߛ�R���.\>��N��v�/<C[>@{�56��Ve�(��Y^��i������@��P�9\Xv�3�v���ɺ����&�"�$�9l���f��g�q���-*\"^X�zL	Nċ˜%?�Φ��Y1�M=?ԟ������t����΂M�/L���������cr�õ
Ӊ��݇󗴥~���M�/R�I�ۣf���Q��ꌉf����Yz6w/�S)]�n*�< }�݇󗴽y���M�1�RN�t���������7��i[%�ُ�0u��
�~N�����`a�*��0��n�o'|�3� �s�nV+���=�@��K���TS�P/j7ʌO�Ob����5�|Σ0�0;�?��bL
)G�F�V�qȈr��<�('ig�g���29W]2��u��6�C�v��j�@^��������� �W���Ilf1(M+N u�p�t*�)N�^�/��Dj{4���,�_��P�D�H+
��
;;�~j��©���N+d��%��[��ͶۍN7�p�����Z";�j�=�'�gЩ�cbk���A����k�۞vn���Ћ^�y�[{Q��tj/�X�6��v/�6{ޗ��l�w�u/�a�&5�I*���8#eIGCyQ�xQ>1�O�f���c�iu^����׽h���*Ἠ{�G�0^41#?��v�,��np��l�أ����yQ�"l�Vc�hjɱ%��ꪞ���j�r�<ȋ��%yQZ9�t/����E3�fO��7�n.�n�jyt=)?Z֝�nb�?�ϴ�꬈��t����斈;H�S�t9�f���B�w~yA�����Z�p� ��fM�����>׹p�w*�)�A��~���<�R?� 0�M�c��_��b�8�h���͚9��j�e�/g��S��'��
GaŅ�~'������V(�j_B}��%3P�>�Z򰭱 �qWf�:v�Þ+���z����)�4���̊O3Pm|G�����b_{�s;\ː�lbM͑�$Ɲ��i��V���ӌ1�6����هUH^�u>nG��˥�ۗ�;7c�Wy����!�H�g��<�<�E������@���sō��^�;�S��nW��h��T�������oͪ�m����4O�?n���������}���W��Or^_~����PK   ��Wtk��  ��  /   images/0732da8e-2e31-48ba-8c11-1e28d7829515.png�yT]�����Cp���;!���k���4��Cpww�w�|3�޼���Z�vu���x���p9ID8<8  ��QJL	  ��@�w��`N���$)��$8z�n���LV@�.� ��P �?�;���|��@�M Ԁ�������Z �қ�v�����* �~� �X����.��9��331� �Uk�?,�r��)��^Ê�~�u��t @d~@�B���v�-U4\4dex��mA�&�F� w[��5�ϝ�]�5u1$v���s�q�'���]��f$%��Ś�TCV�X��ɔ��b"�#&&�s21�Q������Oj���������rc�;�32sss32�0��0�#�=�\����n�v�L���,\,���<ٻ���������L�-�U���_�z� �Ff���X��ڟ�������c�G����I����T������������P�t7����5�s~� �_�/�w�������������h�S�+����i���$l�-�A������/��cb�`ogj��,jogfi��d��q��TeS����G��� 3�_�C����_�F�]����ϩ������z�Q2u��q�S�jg���I��,{����di��������}����?�wĿ���R'S���_����w����{��n�����w�ƿ�"��gu��34�#C��2�>��c��ݡ0��Q������ !�G1aw�i�Q�͈�f���y����m�=F�J�F��a,�Y?<m=�e�1���M_�l�M��(�)�AV���<w⹬-?������&���,ι.t*V������㎲�0o:��pt*��~'��=ƽ��!4h���Y��&<�WO^�Y�Ύ�G%C:Ur$�<9�=����r��}X\[*�^]�wJ���4�u��R�����z\��?p��YyJۈ1����Y�q�E�F�,%i6-5T ��G�~j�J�ht�Z�F=��%3UOYU��)�	�
�p��e4�(ks��(��PNr1����*!���gv�*Fq�
9(h������c�3�3�!�΋���g�~�X��C.WdN ¹Q葸�r��y��L2�	�KQ�����b�J��X��a����F>���e��%�݅�i�T��Ù^�D׽2�� �5P�ع��xɻay]���3�Y��T@*�}3�s��s/p��	��ݢ�L�[�Y�ftuUg�**`B���Z�ƭK�1x��fR1������(��B��#;��Vd���a��9��i����(JZ�9l	���d�;��[��@Y^�(_�Da(�8K*B�x��y��ڨbi(�D��B���F�s�4>�h�?��d�^�v�o��Z_�BKX�w`�ۘ���������:��29+����^|�Z���'��hmRs���dva��7�6I&َ1ud����2���=	B��=W�HT�B����Z&�6�9K�ӣU�O���gCͪ�X��@������`���iG��s��GH>���ӵ���0�P~����]^Y�E<Cŵ���a�VD���M
3ҭ1�}�Rj��V��~�i��k��	�.�vs2$��dT�/�d���x+��Q�ԏ2,�P�@wl���f{޼Z,��:���$��^K�	v��ͱ�L����Da��%*Rx�#	�5�7���*�NL� ��aǧL
~D���E��J�~3CV�Q eh/")�+�10�XV8[�:�4H@R|��%�d[�O ��x��\���ێ����� ��<**R E��*�z@^H�#�����Dǹ�`W��� T�Vn���Y��
�T�闍�tj�o�q�<���U��T������]m�������ut��b��르.�Y%CIaXcǑ�~�����x\P/!c׊k��0���U�l�EƢ6K(TH\k����u��o��`Am�5�&�!rS�6ɨ�By?lܘ?h�d-�$P~�.QZ�S���8����`��o��myQ�-�P�HN�ұ2++t�s�r,:�A<�f�:P�ܰy\_���w���]�PSG)1�掶$�I��|*���gvX,�H+���ah�~s<s����;� pT�(qd���d��N��_�f�fT��%�#0j4��tb�}������^�Sa$����1+G��5&! �b[b܌?����(\Ҭ!��H���7�P��\���Θ��#�=kI9���2T�T�Op��A�SMl8�����?�{CP[��gtu���sś�j�C �H��#�0r�}bS'7� �v�����n]65	����Z�?~�,<}�wK�}�ɝ L��ZE\#��昑���� ��c6��O�p>�xpN�=�6�yn��OMF�n��Ԕ����+ ��$��@O���Yii�-Ϳ��v��Ū���O�&���
����j0/:�M�*4�3��f��m�y`�I����������K��`�dh�9VM�h'H�îg[?�S.�PْL��L���*�2�;�6n�o��#�3��ݨ��J���:��������w7);�˦յ�F�0����xŠ��*s}`θ��A D!a�tY� #����!�U@����oQ<�>�D��b�%;�6�B.+�����j��(Y;p�.S�T�@�pg����8��2�h(��I~�j�R~%�{mJ�Es�^����݈ih^_����� �_#��J(�Y�3�ZM���$��|�8BchXD�h3K�:�L�3�RN�h��9~�, t�D/)�,u�aj�kb�ERv
�,Q��N7��|-D�X@��b�6O��Xm��)��Q���P=M5b=ѱp��Z�C>�1[�a�J����-���r��z��=��W�!����Or�i������b2�Zf��Q�2B`��շγY�(^c��)C�ĳDM���u�/5JcT'MԄ�)�{dϏ7X-8�����w�g3����=��x��"�����<O�#�Qiz m�J?:�~
�to�������ک��V�"�G����̉:�.?�����'���O��T`�k���@�����P�	#����^E��y"�C��5D�33�������\є�����S���@�`�^G��ڏ�n���ӷ˄�3���R�OPw
|�	��CM�c+�����sGJ�5�H) s��C˱B�8#��W�Q'C�$����k1]��(X�l}��!���9>ĩ��@��Q$�U�g_K������Eq�\��@1�fK]f��=?�nc'�­��Ne�X�^�ٲ����h��fPq�yEKZ���LH����=Q����d�\���"� ś�'7O,Q�Uq
����4f�֔ �RH�V���U�]Bz[+M��G�Was�-W�_����!�Klӄf|�!��+��,�����S��gv���1?�e
[(�Y��O�c��D���$��鰁�	!�.ms�fW����b���:=k�O�45v�	�LaJ���!:���̯�K���m��	"-7_�5�D�MP�?䯅+��ʛW���馭�Рx���mT=.YG�v���#�;�s���o�Eڢ��Jr��ll�\	"̄�n��	��'�<�dJ�捃3�Y��<���S��D�;v1�2a]qalh�R�Q�*�6��&�d:\���� �8f��A��+��}��{w����AF ߥO��"�l���C��B�#f���:r��[��ʯ�U+��B����/wM ۭ,��;l=��-z�*h��J$b��#�����֤Hڔ�L2#�*��:���:]�ِ��q]=�Bx�V�e�+S,n��RP3|���W�Oz��*�͑��ٰ)��F���[��U���p�+�p� ���H��{]�*�:�����C${?�ȵ�`,��A/��u}c���������7|J��/�4��>~n��7{s��d�q0d��	�:=5�w☱|���}��:\_qv������Qt-�[����㗗�"^�ː�+w23t���H	n����t�)����B��o�����p�ᚓ��\r�I]����ekE	~��7��֚�����������5~��^��yP��.��w�
������Cd�D�٨�wBV�3ah����jB�*�gF��:��ꦴ#�.5c[�N���=�/m8qV�k��L0�
u:5*9�Y��#>6K�5����-m�F�);���o���Sd������n5USo>���N5�#�4�����S.� �����ҥō���<=��@�GЦ�a�(҆.��'��})t�@��k�-�Z��gx��O9���0F�s���hǄ�"�w.i�E�K���5�iw�V�=wR!ǚ�����51�	� ��ė�}��WM�Y@k�F4�SGQŸ�CI^ح>��EH�ëƱˌ�d�M�}J�Cc#f��v�\\r�,�#<��t��/Z#G%�vM����I����@S��|Z6t��4�}߁-�l��ZT��i�{6��²_C�~m��9g�9=F��Y��o�����&��c�G��t_T'�.P�Lw����=�Ojm\�_����N����zP�೤ڴ茘��O"~�`���sn���{'��#����5�Mto��{��P��r�p �X7-�j�F�l�ZKK)��p@�{�1����[��bjtte%��^���r��<6���r��<��9k��kf�s�yC�^��aOf���Y&.�6iB��t����^->�����h��j&}9��<�t����ԯ�^����������TQ&-^!�������פ�>tIhmA6��˄#!�
��עZ�\�9r�� w���L6��mI�|����h{�#s�#�}/�}I�g���'ѥ��<�����<�@���rS�y���6�ީTU!�~��ڕ=�G�6�fc��G����]�nwn \#a`BJ�ȪweO����hq��b�jR��k�{R!�;�m������6��g`���׍��~�RY��,%F���+d|�?��U,���tT<�hlJ�x�_� �e*����]r��ح�̙[C����^	�����C_�k��K�/h�tqQZ8�H̖O�1���������j��O��&��i5�|ҩ��������Gή�/]nG���}��V�8]��Մc�E���jוj�Te+e��n?<�z��Zw/n׫�(���1��;��������s2����|Y:��x�~{�
����nUf�<��^���=�/���W�^����9]B�xr{I��]>���H�BN����0	4��mTJ�m�Ƚy���C���^Q�*�7,.ѭ�������oj��#��0N(��������kS5m5�N��6J�3>z}���R��^Ϭ,����3|`<&��÷�������A���|̳S�����B�J�=|��'�{��X���dk�ū`^][���T:kl�/�z�(G�V!��S1�����a�]K莵u���[WǗ�<SC�aKIg�r��EV����ŲR�Hƙ5�j�_g��E���2<��x1��#=b):�P �Ҭ�(��_�=֘v��(7rTaJ�F��%K���J�^Z?�\Ҽ�fl$���T���c�fi���E�豔k͕��Ե�K��fG�Ֆ"���s��%+�^
Yӭ�k�������\k�֡�5]c�ʗ�(đ�x)�)lw+���>0"�?��	�\�8m��=��\JW�Y鄩�.�7�F��h���Oz#>6m�95��ʄ�j���Ɯ������C��G��y�L��� �[�sc�Ap�}M I,�~�#���יI0��Xi[/J���U��´�J�8��g�B�ʔ�Ս�%���łD^-�QR��R,JA��T���\S]�X�뾇.��q/�b���Rn%��� �����(��P��S��[Or8*�O=�{���p<CCP�߶p�)#Љ�=Ȥ4����7�e[?jfZ��J��O
�A���2���H!t��3�NЁ�LR�\j��5�4��������B�Z�^���G���tj��4D�Q�E��beXt|3�4J�ϛ�]4VDe=�\2�k����Dqce?x^Zn��#�Wͅ�[���A�O
���
�btP�1$`7<�	���G��QX;?�gy�� F�m��=���O�y���D�����$',��Yt� ("}�?�_pt(���A�
ǒ����]'����)�|;�M2̚�tZPJ��V/5�ޯ���F��Q����7��P��gg�WIPt*,?�m�?3 �iK_"2 %Q:����=z��X^60`?���9��H�o������o��\� A0K
���"X~*�a#Fw�<1w������es��)����^��Լ��P~�qܫr�>�|��5:�W�>	
�a�3�s5���������k>x,X1�:�E�?ݯp,��@�I~��6*M�#L�������CN��F�qw�w�r�Ӝd�/c(������� ���C,h�4���ha�$B����Xw�@Q�ǈ�v���ˁN��gс3"��)}�s����.is� ����<=Q��d���Z�d8��_;7��!��[|�kx/<ŵ��WD��K��uPi���N���wr��M
,sK��&vH���d�OI�-�ܪ=#��P��(N�It�yd�i���8͖�o6���q��&���5\�R^�
�k{����׮pFw�D
��\�5O��!��6���srp<<�ײzzc??���&,�ǴQ���Wq��2;�AT�9��ѿ�R���j0����5w�b�{<�(�}�O�O�+���N���yR�CsY6�x+�����������d�vc�O�/@�Q1w�h����OC���(���[賹�] ^oEL��1�0�0{���LAlw�SVm1�
4��Ά��5]���2�I��O�_��ci��yh�D���&>�����?��#v|r8?��O܇~�1+U�N41�K�Brp��}C��!���i){{���kt��O@g�`+en��؃Cػ� q���)E��]	(���De�)�aC�{
2��Q\HɆΒ���52�$�w���8ۨ��rq��o�㘾b�݊�4���(�|a�ii�j�퓏�f�>���T5��G^-=nd>1QzA#�|��&��%���;=�<t�;֓=o�_�+�a�4f����.N��w����HҜ�P�8�]��T[<�	��H�=
]O��eu�G��2cJ��unsWSh��i�ԏo���/E^G���>/��v�1�Wτ�DN��p.�ю�[�v'Bƿ����p�}W�D�N���9�T�9�v��A+wc�����ש�Y�']�@u߻z�
-ݮ��Ŗ�&�{}���/I����]W�o'So{������׽dΨ���S�Wʇ���V�sd���Z_�(	�L����>ʿM6X/u��G"�c�q�6�}o���L�|~�-��߫������������z�������5�5_��\�!��3)�ٜ�Z�?�w��������z]f�����Z�7�X��V�mk0J���mrêa�����q����W���U�I�^a�NǦ!0$��,b�T=�7�I��F�+�G�Q����cT�1��c��l�n1q�ơ�W�����繦���>�4X��lD��>��u��ц�ǁ��o�������[��8��=u��w%����7D;"&�_��3Yss�ca�5���Z+��f�2��nW��wԻ.���|�Ool��z�|(�W͐�i+�܌��__V��/�#�}�LX�\�F9;/�S@����m�]1qR��_����Ŭ�l�H������ e�m�ҏ��;�|����Uz��t_��T(d�Tc^'M�_��D���~��z[��9��:�q�=���M5��x4���$���$F�L�l��b��$؝γ����5x���]Y��#L�wϋ���|V���Ԫ��u��|�%�؉�aY���R:;N����y��R��'�����J�D��(��N�@uR���{ȅ��*5܁��MO�]4-�1�R�M!4G�'�axv��e� �Gx���K�H�.s�7�K{{!!��l1�f:_c�]�p}F�;�AFur�V����c�'!�f̰������F)ǡШ8\R��\	!�����Zm�>a�'o_��5U�-��&s#̓J�=��K����=�E��ly]�j���i��E��Un�P-��n0k���],��|����D1!�#��e��ϴ�z̭��yx�������N5L	{����
L��v��ۢ� .+2�h�@!�<p�K�~����'D��SED��Я�L>��6�q�C!��20���mWʄ���cuvc~��*#�75CR.��!�~O�=�$/j�u����4F
�O�ߛ��-*"�ߖØ��,��ʎ�C�&�K�2��Q\4ߣp��7�	����ϛ��8�M��E�!$�orQ?��
�2@�3��OPԢ�XM;UK_�(��	%θ������98w[��i��1p {D�H���}��^
�6�.�!!giY�[�ut\I��Irb�߃��Ai��l�Mד[I4M��~�ܐ�O ��������G��Q@�"n��]�A�ؓy� �3�^[[[u�ޏ�cL���ZA8>��7P?���������������&?�N31r �`')����K��@����G����x������|1��3~%�V����]ص�#AX��Q[�&���6YB�^���Q��h������DG�7w�cH\8�z�4�"RA�X��M��S�Fz��mN���sÐ���F�r���?x\2XB`�O4j��]����,��O��Ɩ������ž:�T�}�񒱽Q-��KVU��Lx>\�(Ϡ���󗡚����sQ^��p���p�.i��|�,��'Y#,�5����G�ƞz��8Q�pC9��	cK��LV��Z~ʲ��L�]\)H0��њ�Cؐ�R9����'Ϯ�.���π! v�^����N�7;���PH��{&��p�P�*NN�`)Έ��z~'�q��j�\��w�<����ῳ�.��A���G���m�5���
�G�ئP���xa�0�O5ɱ�<�t�RDۇ`�D�7[>=8��Ӫ
���K
zM���IAl�@���;u�1FJs�Z���>�Crm��*-�<�;$ٰ������#xս�r^S9���xg��u�TH�����{O+��������M��XO� ���b�*U����d$�IpgdѾ�=���n�M�u�w�y�����e��F>�v���1\���	���k�j_���Bb3Đ���c�VA��H�_��:��G��M/
\k�8��͟�
Gg_~^�r�R���{_��M��ǐ�ޣ.Q�]�#4R	���V��.�V�����1��W	����'T(��ǎ��'��R��b��~O�̣�>���B����΁;�3#�[�[Ց	����6���c�+.���}���~pz�!���'C^�s�����'��=��$��(&��W�N��?�k��Ī&���Mѡ@�������^0Nj]n2U|7SK�����N�<�����y��_���A/�O�{ַ�p��|�1�Чl���T��V��;�����;�D�A+�� ��8�ձ�����=������c�!Yxq4�όF���L�wdf��o�g�W=כܠ�ȧ�̈́�P]�el6H��v	.w�5O�Z� ��'�}v�H��w�:�����F����'�N�wb?�[����Q�>�xZPl�X����p���2�$zr��S �����)�V��RI3C(2�c�wz�����D�|��bZMϧq���Ӯ���*�֎�n>���B�j df���H6�,�穊��,��;���^�� {�P����-\�P�UJ:ԌREn�E���
��wpԌ�Ũ#�XZ��6O�xf��?�&n�h�}���Q2XL�O-�Prw�8�dn&$V$�Wf�v1��a��NH�ܐE/UI(�*E��g� � �y�MBR��hI�x��S��'�?Z���_˂��l�´y&R	J,�[	�j��׮a�g|�����.SV��#>X��*j^�Iޛ��ݲ���)%�yz��'���{i՟�v<�W^e�|�_���Y�2/�X�����t��~�����*3e���7W�05�E��j�{L���#ɀR��"l�հEM��1�����F�@���d�ޅd07�$��5�;30k�&!�U��L?b��5�X��[̱�==0 ��͋�S^㠐j��!ah�X���R�Qo�D���Š������F���[Ή�"�O0m�d]��"�zƑ֝�E���6a�NH7FwT�bA#K���t� `��qf���h��LU�=>��jP�֊h���JNG#� ='��������!�I�(o�֨��o�h�=qIN��JI�� }^l��� ɮ�l�~���#�?���i�q@�Y����D�4Z�}�:^��c���C�ݭ�쉦��m+�@���,�U�15�d�9�B��o)��>�p�K��$ģ՟�
m��%G 2ϑ�w)Eߝ0ɸj����M��xAU*��UbA#�[�.�����u($���R�U4Z��X�1��^?z9�e-��i��ž�Yh��@S�m���,�W���a6#9���P�D��Ag	(��f^��*0��-�#��7�N��wa.��>7{F͊�Q��2��/�d`��JF�7I#� �0��i��L��g7�Sƀt���|�u����9�~���E�\%�4������S.ڪ�ܛ����1'J	U��e���!�ǹ�-�;H㊵�SS~�A�)PZШ�1z�b�/ưk	��8�pfb�}H�rҿs�=�ά�|�=���+%>���� C؄q�yW��$��n�@��u���=��(�習��\�d�hJ�C���+(��v9���&��0m���$���*��+���}W�=�x
��"�7hٺ�ac|��N�3;s�0~rr���alN�1�YD�)�[ﹼ/\H1F��ݍ��(��/X��%���vJ�%�k`5���u�sv���/4���!��,P������O#&�lA�5���Л��4 uՍ$�L?(L�m��T���ST���Y���Z�����H`��|O�cg|�����X�h�)�c.֙���mNdT>j����@��PI��I��B~g�����0�@�9�>��ˇ˝6�_J��u��Hx�8��}����0S���S� ���~4>�b��ۉ���Ǌ��i��+F��E�g����|��)�~ȁw�kȄ|�'�M�y)4aI9�����Ӓ���<grj�{=Y9$�]/,e�ѭ��w>Q�#ՠ=!�b'�ȑY�� �O�n�E��8��
q�[��ӊN����៯ES��p���SFDU:-`웵,�%&
$�v?�?BP�!��y�%]L�"���rG� �hdl'nQ��01�П=U8Q�x0��}���'8���@���0ڶ^���*�a����\e^�ږǣ����z��!�� X��8(�T �̩�?�� �$�Mo����v���28��z__�%r��V̳}_=�u-��h�dP���2:���\F�8l"9�.��[��}��u)	YVR��@�w��73�����~3��q9?��i��G:>��F2v�!�}blV��������<h]��|�F��@��Mٱ��*�������|��}V4�%|&8�F-=ܥ���V�V&ݭ�a�`���	���;��%\�+ <\=N�Vk��I����w��R:o
Ou�ŃKbZa�f|f	E�r�9���gg�����g�g�J0a�R<i1B5v(C�=x�ҿ_��c6W&�^o�%P���zF�
�\�/z��_#I��.�s�O���2�
7�`dkZ6���������\�}9:��g�˯�Џ���Y!�(���&�蹿8�Bn��/?1v@H�D`���l��n� �n7�xɘs�F��ű�` t5��K��w��^�}G�c�^F�_F�;/ �����,�ſ�;6
�>�.�b���O������N��DP����Vq]`q���?����$�75�@�o����f���D�L3�� ��/�nN¡����2��3��A�jj(ј
B����:������T/�'��J[�z���e�j���ϗ}�j�.����_�.ti(�0@��&c��(�Y�0P��h t�(��6pH��'.M���:	�u��AL��/'���3�oOK`�
b�����ز�V�A��TVa�a!
Az�'�k,���{��`Q���r�%I!S�VP�|���S�o/M���ѷ�g����.+�2���]n�E1K3G��?��X�F�H�Q�9��"/ɫ�wV�+�1-�P�dX���k�<��wlj�0l�K��}ۚᴀ�5�-3�*!�!E������ǈC��.+�Fjn���0� ��C�d`j��YF4�q�uG����9�ko�
��N',��*�f�I�GFP�!_��.�5��Q�ݵ��,�F�?��FT;'Nl��&vr,�NC>|�94�[hv��J��؃����O8�w83_I� R[��3;Fk�?ٞz��h�"�9_�f��Y,�Ba" �rƖqr���0�R烞�ZQ&�M��~Sg>�J��`g���.���Pmd2�����&�X!�i�F8:��.�v���lRl�"$5j���"���"��F����{.����Z��F�x"(�D}��m=?4v>)���K��rHs�{v�{�X�	�Mئ��) $A4��GF�=d�|̼mp�0Z�(�

���6�#�5@�u$JONuWpi�\�H�碏.C�\�u0m�h� �h�>v�]�_K�"5�*𗌠A(�%�؈��{F�]�U��f��dzw�J�4�)��'9^꼳�A��tw����@w!4�N-����w"z�4�o(��V���јW�%�d�.]G��b��J��p^ ��>#1W�~_߰�fÛ��1K�O1�1�F�����A���V�m`�|k� �,�F��M�[�o�8L@ �	�a2��MX��h<Vs�j���6����v~�tN� ��:��q�-����L��C�_OM�3s����P'�h[I�C8"{A��l�Fq^4+��qw��P夀t!�>��J��M�\��Χ25�������,�X_��H���
��;���0��4����.�����y5a,�	R����H�b�\IFaF�un���cV�5�8iQUzy2��u�꧗�8'W�0�hT�܈�J�P*�f�bO���;�����BT�`�&z����U^����G�X�'�x9��""�,�g�2(��=���T/�~?�sD��]�ޠ��bH%\��J�jr&�����am��Ҹ3��#�RR�4GOJ�dH`�^'+l������~��'�痢����1z
�q�vP��v��D�E
d�(��t�X
#�!�����s�r��K�����a���Q�d�K`����uu>��&��i�0�f�`
]��=2��#�{ v� ]�E���j��'�B�s�mM��&v]�j���f�iZ�$��}N!��S�o�0
B���������|w�<x2ˉ�w�/H;���ze�m�_p�8��S�!8�}n��.L.�p�s��Qi�E-p�F9`�49H��r45Be>��qg9�=�U����\(��6�/�N�X�C<�R%%`���T+V�P�}9�|�ꩱ�]���(4�X���Sd��XZ��xծ��p���^&m��!�dc�0����A������{c�+
�D�fv�GLsB�6b��oXx��9�����"a��z)Dz�����Uf4_k��Qr�@!�A��W^�u����|%�.�X:��v�{�����33�����S�&�,	�ٞ`1�鞜��P���]���=[P%��B�"��k��+��sq�rēs�v}V��)��:�w�d_�ioP¦d�^���FH0
�e߇u{�qWvO}���%"5�W��/�Z.^�@/��v�u��1�����%�
�Q�`�m1E�$ۉ���5|t��ТKZM��C��WӸ�n�����!�q��S�/��;�W���ٵg�ŽؘvP��҂e�31.`��	0!�����XYҢr
���9X'��CAN�8�q�^������j��h[\+1{$�d��'�ϓ�*9�Ąb��l��pZ�j�XM�r�2�l��������^`����aY��H�W䪜�*I�����
�'2�ot7�ٺ�'HJO�K�|�E�?*�z�����eG%���xr��=Q�f�5�!�t�"$��s�蔦"0\e�/��?Cg9���+"|B}�M�\���������'����o-����>���Ot��f�]𹂯c 1q5Q���ad�Y��賙#�f�������O[2�	\lA04O^�29V�B����8eC�Đ�D�[%Lf���L�+Y�(z��Q���bi]����w�tn�z�޷k9�y�����A/n���+YFr�{�3ݚ�f��y?�#E4����8�h�����(�<U��9;���+)�<9L����e�%��^r��1d0�q=$�K
��@�K%O�*�9�`Ff�0�`��7��T�>'�T'��#Z6�[��m�q�m��(�FD��P�*B�)�� �+��",��y��{��T��`l=?�䨇Al$PdMzA�p��i��R�d)AD�`Z��V�=�Z�������+�8|C�|���Us�it�G�챮ߑM٣��<�HF5���|��)���塕Y�Ы���7��)E�{>�o�-�6��x>��69���M⨖�Պ�����`�K������O�=��*��}\��a>>0���Z��|*U^7�=ݞDѕ@������ˆC�_&d�e+!��暞�}�Z��v�j,�D��ޗDzw��@3*�U�h���{�����+ƒi<����o�gh�س Dζ�����C�@�C��x5�w��Z|xƇ7�� MF��(�Օ:1�G�)�S<5hQ��I�� Վ���奄��+pP�4#S#��HÄ��i	!&�}V�X{��a Ks_��롤�Q�WAq��f��`ю���"��!�2��1��.���+�b�\Wj���4x��8i�6�U�/�P[#��!n:��R��bhaĀ��@�P6�������^AZL�[����1�פ��������ZN�
��9\$P�����φ��*��{̺L�=�t{�O�}l�`F#	��d]����z�^�`�]�K�p��ؕ��P�(mn�]+��84�`XN
y?gC�ZP�q���p8HdD\��G��K��6d�Z����\b��-��D��vQ��GLq�H���#%�u%p�g���ڞw�޾	���	/�4������G@k°��y�s=6A��k ��lt�����Ic�}��4R���=��d�]d2{�$�-�+%�լ�8��[�$�u��+5x^��mO�hUo���8��s�9L�������rz�:�H���-s�8��v��p
d���'x��{�̻�=X>Z�t�ѐL��N���9�q��+S�]}s�9(��T�U�85Y�vq;ʵ�B��.�"4��q"��I"�E�ۦ�W������)�
G�����!������
<}��&H�ѕ�ERsEUq�� ��}��m?�����R��vb�߀���YR:��9���"�ѱ��p].�*����ѝ+,��8���f�=d���z�ؕԒ�Ki1�� 1��������<s!u���;���Fi]+B1��=j�-֣g,$�7���S�RsއJ��Z��O�l(��"��H�/�x�L���
�6���\7��EǄ:��!P�gdk�� ��t��V+�Q�QYT�͚0�K�|����c�<���d��z\�Io�8���4�L�[���e'��|�3[�Q��;��J��o�|eQ�0�B@*G��c� �̖��:����` 	w�yoaCO�xޜe*�$�bl���h����������� VR��&�S���H��%b�|��  l��?}Sæ?�kn4���6���8}T�̾�,��Y��*�EW�~U5B�K.X/S(%S*�]�k�,��z@v�QX7i'��'�`��t��M�S�F=r	ti�>&�+:�J��L�X�v'BAe8��2����>憐�&Ҫ�κ�cw��-�N�Z@�}�2�~/WLGc�|^��_i�'l:,[} �?=�ƛN�A���c+T�\n��W8��*<`����+�����| ���>[�j3����uE�;�����G��%�6s>O��\wy"���ʨ�2hP�Sy���Qb4C"*+X��$@ۿ��_�买�\� 	j`��,#�%m��&��P�2²���e7�H$(�J�}��_�j��c��V���~�_�[�n1ega�t�J���h{Y��b ҉�GT�0\ ���$��/uF�4�6KS(;�z M۠F���W�.�[1 �B�p�� ���Q��@�Wr�M0Â2��$(;� ��K���D4N`7x��U7�(���%r 9A����G�VID��ӿ<�z�'��,2)�AP�I��-�=���J� SC��u��k��n�r�>ݖ�«ʛ�k
eQ �W�)L�����R�S���U{	�qX���Ah�<��XG�v��<��SAB�$�N|@��!h�U��  @ IDATէ^C�l� �x���A��l
j�D�����C��qr� �HP���m'W�)��B�N����R���"���+q}*m����1��@�0:�6�\"�l��D(b��q�D}*���л�m���� #��2�f^m].J�t��D&���P�HM��]�`�NA���=���i��i���k*�Z�MT[�b�&w���!N����W-;��Y�BP�:4����j�>�U� Y�2�9N�^���M��'�<N�0P>Y7,�c�,��;�t&�t��Ut�:�t�B�D�@0�B�1n{�8��u��.N�)��t�B	A��U�.Z�P7�B�Q�d�Sk�-��]$����\��8)
l���Ť���Ȳ`1$�(��K� �W!��`C0��fFO@k$]=E�%c\�A��W����?
�e�`Q4����DK��Җ���>5�H-e�:�=���ȷM׊,Z�5n	 �:Td�3cw"hM�H	�:9R�5hgn���E����5 �S�h�Y��~w���h��$j������*�����s@= �2�"4eh�&�O��J[*1e4�Ҥ�R.NM%B��?
�c1�׊ �y��c�m-�0���霆$m�A��3���I:0<QEh#��}����������(~��Ȱ-ks�T�B�l�4r@=4�2�� ���!E�na�zKn�Wn
������`"t�6)g]�[P�-d,ݖ��r >�sGg��[�"�V����%��%@E\_�`#� �j�c �r��T�D��)ޢMP�Gy-���H%Q
b�4QIQH��>-f��6�"'Ey�SY�+�z�E���j�-9P�C��k�R�1��P�=�����h�R�""6N�WP�"n ��
�O(�\}���KS\�%�( ��A4cD�M�j޾�5�q�؍�BS��] �P+��>rL8@/�_�e�*�)�}�.�' 0�Z�^_ݸ+3��a_��1< taPQ^��o��H�z�M�1�˥Җt]��t���'�Ͳ��պ47�^�HW��?�A䬌rE\�]EB� c���Z(B���ET T<,B}� �fj-<5�V���6���}u��t��
+{������q��8��>w[��+����"q�l�U'�Ǭ��*�
�h}�م��.�90=\	�AYeϕR����娇��G<�!\o�P%q�?���rѩJ�n���ߨ�)�[�'��q�g��8ݸ[�8=������U�uC��ȉ�
O��z��{
=��*�Lŗ��vZ��Z�Ʌ�e�Wρ'�D���bUϢ�2���������ګ����@%�i����aY�#���%^=&�D�K���t�>�t�j\s�35�}Uӭ��*�\�M��̅s�Bڐe�b�Oܴ�kP꫍��6�[=�L��~{S鮱��q��(ڊٕ9�N&�`���WAmA��!Z�(�q���,0�����E�%7�"54����~JR�U�SX3��/O}��G��Zg��Մ}=�$
ھ|�r��'���HL��R�r�#��6^C\�z�p�1��̭�\�(I�1j��vg#��?,8&&:��!���H��Z����[�Q�����w7��td�=�w0��LskQ�����������^=b��ݪ�P8�̍<���W3*O}a3����s�F��tt�vkp\�I� e,R_P�4z"AL��AE�6��	�1���3�bBCN�z���@�sП��:l`��+0|� ����+ds|0�'��f#�����A���'J!mV��P�@QJ���������|�I�Au�)��3Ȩ�|�r�!�<������)+��I��N�n���.:��"�NS~�f�Ӌ�)n�����riP���ǔK��(�'�9��K=PN�#���ȱ��^7�$2J\�b�}4A%���$������OQ2G̛<tD��X�9 �9�2�`��z�n���jw�WV���G�1�K�M3��p���H�$�k��q&��RL� �nH:n[�yx&�-�SQ6D�+�zZ~�:��m�aI%�U4E+Τ���E2�U)�4K�;�O���3�nsVY=��Uh�b4��	�/׃P/��2�qB��~��d�Wf!��R�7�΄��~f_&�j�0�������Z��B�R�L1r�r��7�K↉�#�-.P*U��Q�i��"�|�*�W��ڒmj�Z��d��]~e]��;����L��(Lg�Q�Q���h1� ?3�I�����7Y���IGh8�"2v<UGF�I3U��m�f�O���Ƭ�z�F�S1�F��j6��
�L �.�ƍ�Q�Z���6�k�x1'w��[M.�CF)Ⱥ����R��v�^ذ�\�n��H]n�~\�H5;He��uR�Z�m��]��JQQU�pԃ���ۈ��Fs�|!��d�V��	�j�ޑ�n�Fes��Z���=~J��jt[�r&�Te�9$���n�=W���PW��v;(m\{������KW;�.�d�*ׄ��!���3[�>{i뒨�$W���v��2�USW����K$��֏����?iܹ�J)���ߩ7���x���T>Lm�eΗ��fԭ5�}z��è�L�76�[���r��gfR�l���hAo-�ߑ�٥R�!�����<Ƨ+L�
ѽf��g"d܀���.��7k�{��Wæ�9�^/�Ozw�N�K�^�[�c�:kk�8s?dx�u�(�f�*&�X�\�H�I��*������R�]kdӨL&;�nvv~���/���S�p��w�Ώ���y�>��>JG�������X-�+>�p�bH�S���+	�<+Qj"�$p��c��(����?�������?��/��f6Uɖ+�o����g/Ԫ�|����nP�e��xP�҇{�?�s���n���<:_�Wr�L���S	xk���K���Sa<"Q]K�$��t�
g���o�k�7
Y4M�A�Z[��[�0��)jo��'1�M�n��o'���M(��L%݉�X��b
M�ҙ�*�n�FD�kn��,�Y�<�K�dB���Z/}������SW,�_(�A�P�u�]����?��������S�\>ӡE�:`)m�W$���cO$%yt�΅T�k����i\��>J�ڙ�Zm?���t"�A1j:��ފ�A�m���zm{��s�5|�&��n���2~�L��dA�*�@����,�.�	�".���f��1��̅��:á��sX~�D�/j�j�t'-�ħj�Fʬ1�.~��
��N��'&�@��IC\*�EA��z������&�2%�2�n���v�P
�-Ə�J9����V��k���fuc3&����8��1�Vdҿ"9�Q���\��zh��ZZ�3��ݿ�h�ڵR��C)R�J�1�f�T>�e���l)j7�L�k�B�{���0R"��b���<��d
2$+#�yq�����ƀ�w`\5�#͒.��L6�d��DR��n .O����P;I�����!r��U�J.�L��L���	l�R��[�b~#k�fm� Q(6��b���Q���fO��t��N��R.��N���b��j:j�ӝG�n�z�"�ɞ)N�Y���~���?�b�!��*O: h�yX���f;��V���Ǎփf��_ku��J�SG({-�?��k�rZF��F��IF��b���tD	B$"�aj.��JT�M	����'���&��������Ԅt��X����=�@L6CL�Py�,G6Cd�#��y��f�_�c�
�W.�E�@BQ�I��Hw�A��S�.��V�xн�m�a�ɤp�N����I,��n=�熛B�J��{�R��_?-�>��=H[�j��]x�˶��2oH�J��6.~O�bC�q�e���Z�ҸML'�L*Wγ���'�P\� =�R_Q�� 7+S!�L"���Ujї��V,#������9R�6�@I)�Q�($z����s�~�F�(ì�qbnēb�nZ�F�������C]Ν�ʺn6�c��Q���A���m�"�K�����B��)4�,��ґ��U	��m�6k��CDU��S�{ҙ��0<�X&��EA!b�F��|28ȏ�Qqݙ<g:2uE3���ɓ�^���2�	F�p��/9�%��`@�
9�]Ȩ�ԏ�z�*d�6*�3�����2��G�²����'*���T\�"��H	� �t��6Uwz,^׋�,.b�It��ԅ!��7���b�����ԻQ���J6m�������S����"��VM1�����0�OG�('SLΏ�a�&#R2� ��W�jԳr߯^��n���e`!Γ�Ʊ2�#��8�� �cqp�Pp�q��K�E�"�D�a������.�xB�J����M�T�o�m.<O�zRD�3a� c�j�f��:4�>�����%C��~�Nگ��iqԄ�I6H��k,Q�3�W�.t�J��6h�Ճ���#�xLf3��^wX,�K���S֮��M���݈���B�+�O����2eX�a�f�F�(d��n��e]Q��0v҅L'^$�[\e��j[� ��B2g7��b��� ň�B��"�2�q2��e��و�t��/1�3�`��}}t]�e�@Fw���#J�3��6��skklV�0��O���'���;�"�N��)�s�R-�h�XZ��Rӱ��A�U��lW_=�M�d���b���T$j��^Hu�#�n�̙��"N��'ޔȌh�>8J(�1���!��b���M�-�LP��i�����
<4A��r�(�*��F������h�96%�;B���&
B"��x�2�N�.A(Sv�^1_@����D	� �1ߐ_I�:{�b��+no��<D�B3�n�*���'8
Ccԯ�z0����+"��")6�Pu�G3g���(��9�<�xt�b��[��3��u<�bQO|�f_ E *�pwe�4�Z�0�Z�!'bf$kFj7��c"2e��n��p���0�%�I��5� ����	�;�Ҥ�[�+��0N��[r�E~�� 	��aE':feƝ{$�щn���2�B-1+g�+W�>��PaM,�Y<��$�'�2���E7n� �OH�U�|�����%��H>�ٹ���d��X�`ߊ�Wr�����Z�͚M!bi6/=�j41�zC�c�(U��@��t�hx� C
��bU�Cήj9˔]�Y�����Ϭ_ި�>����fX*�&��P�W1
}`Rk<+�� ����?�� Y*F2-a�o�9��v�& e�L�嬫�L$	��ʈ��f�4IGx�!��'cL�	�q�@�H�9I��n�\�|���� ���P��DIL��Q�s�����kk�|��9�6���TnL��$��{�uN�����#k[� ��z0��3�����ʗ9D�ߨ���v�|7*!�,�B)*1,���	?�6�!�H�ȦJ��d����<u��?/�i����O���'s���v"Z�٭�ǭ�H֠�ҠZݗ��v�g��7Q	�$q�Q��:IEK����!�QZ���d��@�Tb4Ȑ%/�h�Ī�YM�pM?Ҡn�������_o|�˯_��y�B�ݑ�;�`�"F�D�dW��ci�\hX�a� 3�3x#�fT�� V`�i��F�Ĝ��@Ȁ���?�r/�?�;�'g�U���"\zV����3�Q'ԁRf���Gj[�M��Ȃ�2�©�l�����f;EL��`�}F=���v��&_�H]��X][h�( ��!͗�G���_��j���Qv�Uݯ�ഋ��wo�*˭f�����T��~�Lv�b"#u? �Ȝl "�ȷ���L1Af]�̘�<��8�.���l9�������@#�<P0�f -3r�\f�K(�<���m�I �W��PXBC�����YFۥ�	P��rf3��ђ�59�e�Q���Ҫ}D��g��nK�n�
�G�\���z&X�����L>���j��"4!02,�A���?:͚�̿Y$��6�"�v�.�E^�}bV�x.�/�&��@�c��̳��JY���F��	�FK�/�窍y�~b.��A���j�� ��"��3�.gd�l�ޱ$�_��OC��"��!���"��2�v��V��u���M4� �Tj��"&Kc�1����d�e ������'���n�8�e�'t�?�m��x��.�5z�$V�Ȓ���'���X�'0X3�"z(��U��e 750�3�E^�-dC2�5�Ʊo�T$��w{-��A�g��@��F��PEul�%�
���4O����6���Gϯ�뱉ӎ2��5у^���+*������@k�.� 3USH̫rCć��r�6��p*�Î
�5בIG}�ŉ�t)Ğ�A��8R()& *%��y�mu$�/:��X������www����7^�u�
#�f���+����@d�]�� �"7!�N%��0�J0Q:�AL�w�p��D��Ƿ���k�.����Z��:�lm�?���"`�8��A+يG��Em��	J�2a��2Dh�
}���G���wu*��v�t~�S,����[�̗JXm�r���;��!A���D,F��?:ke�	�/Bs�y)��*�о.h�~�;۩�uf',�2]�
�)F{V����� �?VMQ8Y����fnć�5�"�']A0��~���C�Yl��T!�E!ۑay�T�V�1��}$��gL�bAb�4�Ɯ
i�[r!�x��d�Ý�I���0��j�eMRd��aԅ ���80ꉗ�����Oϋ�-��G���K#�U"�(q��\ �Hhȑ-�~��"V�X;8) 6,��Z�ݮ]�:�����1U�̺a��^�R&�����;�w���YYn�|�Q�n��W=�D�O�,�ɢ��Ǻy�����+/��һﾋ�U�k�+f,�R�(��f���f��c����"ԣ�j�	0��稣1k��G�b4�"�UeY�>�!f1�u�E������� �b+DSȓ���3�,���*��8��[��
�����iH�!DPą�z�����Q�R���c�"�W��3&���"p�I���L�=Wd_LA������P���9�.���"W��i4�o~���!�.֦�b�EM���nh����q��Fr�Cbb5�i2�u�	�(�<,��L [�1�Q�{�U��S��֚�Q	B?N�W$BC��0�c"`���<6�+sfP�ʔYOw�|\(�Qpǿ�+�:�#׽�L����]n瑭t����3��K�Ж�/B�_ǚ �|Z�Ɗ��	�d#�r8��S��6��Ç�k��TP.�PdfW(�X;D_|C�+�G��*r��n����>=Ks�h���\QxQ|�,�j�F�������B=�Y��L7Fd7���dI�3��R,~.����Uߚ�I��C2�|�[�@| �^1������g_�C����	���%[�f[Po��+�Q�&'9�n�u���v�|��^.W��L�U�59{��Rh{��r�E���hH�N�29��g��?6��P"�V��Z$í\��G_|Y�0�$4����٨�è,��>�1("����{���� ^� H�F`���J,�a|��?�A��D*|^� �,�źS�3h3��T#j6Ru�-F�򅌨W�t[|�K,��2�}��N�L�Yo����n��x��[o�����08Ų^�`A�: M��fS�J�L͹8�^�e+e!�� �B���e'�g,��;��YA��Q��dK�Uvm��m1|f�?�.�H�:�H6�e��Sg�N|�fd��hϟ�e���ΰ��B�g�D1�[3���řf�3{�q����)��|/k2�t�pI6@��0�.���'D@(���k����0I�|`����ŒZ	�R��_+�xŎ>��VHC0Dxb�
���S���÷���9��N����2��.$& �Sd"�Y�Ӡ���P.�܄ה_+p�a�Kmqi��Px��9E%s~*���lM��|��\yoo��,YP��AJ%�avQ��=�}�]Β��E7�F`�F�0���h(h H��pA\89������*vcq�l��ƃ�������i7�d�0���<�3� Ks�>TB�#Vd2pڵ HrM7��L���5rsIa�ë���<��Ƞ��Z�7�c�)Ngawo��'Ԃ9b��2�h���'r�����(����=x��0�[崨T(Pe�cQf`�o8L8o|��>s�xuIL�����с��Y�';�<ҧ���Q�d7� �4U[�p�8����~E�3�y'f�x ���"�4�(���s����H)f��D�j�O0o���	gi�$�A��On�c#��\�E\>�3�K2���AW�Xa��k,�p�P!��_Q�\ܐ�+.\"��[�.C�P��:=g��E�IQ9æ
?N AE��nq����YuoJ��J���t�?��Q��ϙ3g
.x��HG��E�U�o=�c�@f�(" ���N�:�|�V&!`H� �Nr�EW9n�_��g���E�,�"��R�l�����v�N��>�lN��Ĥ�θ�X�1��cxY�e�P�=De����q��d��V�����7/F��|%�7�.N���셛�Ivȯ�ߌ�b=䈘�O����e�>I�Ѹ���4��:MR�f�Nt���<�e`5VS=TdU�h�v)�ָ'r��D�{Y\����\�Y��3��eҺ�/�n�>`���lf�E�٬ "d?���y��	��J�E�fu�D� 3d�$�T�b��3���ʑ+.����-G2)�����r��i_}�2�7^���UH��;��.D39��b�B��/��C-���]3Zq��UT�,� ��V!UTd���T�A��v3OtBN�.�n(��$���"��|�:�2z���MTH�o6�e���ѽ@�)�K�'�d�d�X>G��U�D����0�M��MX��Њ�&����S���Z�����2�TcȤ��/�wf�Q��/���D��F����15�$�*�i��ҁL~8?��I2>a���+�}��YJ=jUk���q,���WJd�V1�j�C{JCFG�0�+�p0Fr�?&#-b���A�Tz��,�RF��Iq��V~uMV�� �I�_>�mw�_]�6D�8q��d9�8F�f�3\ـ����9��:��ɜI�dT-CMX�"G�!{R�ÓO�X]
R�@)6��lq8_B�z�61��c>�2��Aw� �$˰�[$�ڈW�rQ/GWDQ�
�I}�\,�.}2�K��R�O�޻���W8s0x$*}XPJ�z�a��\�CiY5�m���	f��P!��8�K\ב�û��A:ݚ�t�}�F��#I8*ئf�,���S�S���\c�E	�3m4f�!��)Ey�n�촚m��@#�Ԁ
�IH7������,�u��J���f�T��*k��s�>�j�F�/F�Y�[���)c�D]��'�C@1�5���c�f��]+r���+����M_��j��:�j4��a3Þ�hR�|Y�d<���Pf���S�4?y�	a��-=��/�C�|��=*���k{�*�[gw��fU~֩�;l-�J+���5٫G������da	ݐ���k� ��Cm�
ߕW9D�����w��-������q�#
�mʕvA�k~���Kj�hrD���f0�%�r<�?E�$Zc���B��$bC�D�a��ދ{R�f�b���1�����G�Ͳ������F��
�����=��\��B���
�e�|h��Ň�|(�˄�Au�2rY|/4���9��7��XY�o`E�PE>�
tT����(�wf~�@\~��|k�Z����[�5�¨��R%ڭR��ឮ|��zd1��������ˉz�*���G~�z�����Jl��nX��n�K�Vt�*��6j#��|�E�u�mh2N��uؔ	��W�JqSEXn߹�R0?b����X#L����W*�ǻ{�ﳕQ��)��?�:w~�T�{��]�[�ؐt�����s�>�pyi����~{-S����M�'�P�%"����zS?'o�	�w?���Jş��O>������޻y�����W��������[��۟�����R*�]�����݇A.��η����=ھ��{���3ΆDE�jY�y��eV���2GO��1h��a� ݬ�R���ܹsl�P�!�z�#��z������/�Y}�v2.�SNv���a�h��qb��V_[�r���J���ݻ��_��������{��f!�m@��
��ݻ/���������n��a�z��k���u���bu����k4��5EV��L=����_hb���KK�3��(���;���kս|����1���N�)�����>�~�{�V�֝�7o�a��Ƈ���������n��r��g^y��{���T�Ł3�.,q��B��D�;a=��G�%p	(18�a%�2��CF��� �Y�D'�8^��#�\���z��#����fV6X�K������'�J�Q�z����Z��̕�O>�(T���W[�Q0�mJ�fY���U��Lg/���w.�+�p�����n���I�R�_l��Ŝ�|aK��H�Wm�2ܢ��8w�TZ�~��N�6�]j��݇��z�Re��_����>R���ō�D�Q'�/63��j}�ޮ?���ݍ[�t�om�M>��"�r��x�0���ji����|�Ǟ��	*�t��4�fP���X�V�-0{er͛�3#w[-�3C��Hd�:�c�����L�V��V�sl�����-4��J��(,��v�Hl1])6�k�Qgs��z��pg�|n3×�a���z�ɜE��c�fYI�T1C�c���*��t��o-�rm]���s����F��:����[�fg���rr�+i�z��V�T�4���>��Gfvv6>�I�����sg��U�4��kjW��`IN�n�]��Xo'W�W�m������-�kF܂�E��^R��6N61z��و�KE�I$�-<�����L~$��:�kdFn��U�U�N�3c��cFdY�/6	�#\9��!n����			1X �`$����lal۽/յef,����_fTT.�U�V;�&;��{/��������'�)��B8�r����}׈Z��W�^�O�A�V�l�g��(�+�L��<�j�`@'��s�Mt��K5�Yj��6u�,;�X�F�G+n��6́TK��vև3�Ю �"r��m�S+{��޸���b���sg��7b��͏��/���o�{O��'�Ƀ�����}���G����"�/�
b��rA�y�����i5�#.�������ϥ���O �
�p�-�R���G�r��ҳ�)o\:4��W<*���rH��N10_��U�5����ag\�F�qus��j��(x�̈́k�%��1�|F���8���lmo<:���P�M�PG��D1�0��a�6�G�>�9Qp4���gU��ؾ|�̕Z�^��p,��AX.��\1L�B�� �1�����������ݪ���������j�J~v#�4.A��D�v��Ӯ��J�1	fJ��:����4���>1J�Ua�Ks��D.}�ynI��B[�N�5�=�����au�q�0��}{����g=l��r6�9�8	���"��oP8`�F�NP��f���+�~t1{�3|*s�6�x2�ۀ_�)�J�Z󑡷Q[o]�~m��V+�u�v��d��N��h?�@,O<��ȑQ�ß�1�A�a0��[�-������ݻ��'R�fGp�a)��1QڕyAЕ�}��V�Bu)��܌��7�ڜ�y���7����>0$ݥc���\o�;��^�Nu���<w��B�q���a< �Z�'~�
D����|�u�#��e:����´�n�}�5�d�"�Xd��y�~����?�4�qf��e�����pS��9�>��K���9� �ջ!.m]^��s���k�	�E��bi;��_%�9+#�CN z`�Uo7;���^���_��/ɻw��n����VI��<��!tP���|Z��2����GA/ 0`����V6���iVS��J��mJ�h�"]�b��t#f��A�⪡���S�Q�������(�� A����53,LD�G�WF�pac��{��?W�Κ��m 4!W�ی�נIm�e�|z�L����{���:�F1[h�GT%S��eM��1�Q�O������07�O�3��΃��r�����f[�*��H`ap���To��>f,�����kGB�Rvm�-|������t>:��!J�q��i�� `K�&�N d�v�[,���3�gj	�43�zaS�_�(�i�>z���03�:Z�doO'�c�?��R΢<��q����r��bPF@�96�����7���[wƽnΤT(�s���X�c[����Di����N>
���:���h����r4AO.7,���q�F��p�����!�����K�p���]�Ə<�ys-�f.["�|�` ׈�F��s�y~�R��;]h7���'�n���1>9�7@�0�-4���0P�Ň�i�b�P"�7�f�V�^$"z�tj	s��[���h�U�����^�U�6�:�B+Z�^L�#pL��X��g����F��x�R�w��77��6�o�4~���.�>�|��	?Ī��~H��õ�-�|�[�7��a_�$7�l|�b�s8
l�B ���O̺4��*�	�p���~����e�����nݺT�C:J���ۋ���^�����O�m���o�q�s���^��F��*M���0��a��/�h��f� 8j�;%�KtP��� ����H��s2�˚A�%+� �n��"l��赻���fGt�����:K'BO��^��@%UXpD)��7$Vb�@��>LQ�
������������?|mܨ��[��ݽӮ��a�1b+�2�έ"�����ج\�P~�d����ׯ]ER�*x�G�kMR0��A.93�@"m�6�y��ۍ����g��vo�1V�ۓ��XH���eݐ���rYg�e?�����On�՟�1���~\	ⷮ�M��@��T*�A��8&�!`��XF��8�a��9sI��M��#t}����`�en��t^C,w��m�H�K׬$g����2<�5�Ѥ��s� �
7�(�K�=�onf�}��A��d�f��l:����C����{��=ܫ����������rP$F���㸢��m
b�F#�*�YB���D�
�.}��ԇ�݃�����/'�21�w,ma���S� >�`����$��pJ�_�a��bKBb���K2/p�G<�=�.,%�;`	Ě�R�����=��!C�8��y6<���+���B��8� �oaJ�rY�Ѣ|�RC���Rˆ�=�N`�a��ˠ.��Ӵ
�� �~�"KЃz%�s�I���� ��(��A�+(�N:�8��kX
|�KJI`w�{�(|���g�0H  �x����V�QsK���\�{p��Ne�F<y����:�[(!���٣6��<)\RJ���pΒ�y �A���~��X�)��(�� �׆�a�qh0i�ol"K�w�	�ƶ����O+�.ĭ�4�5pa�5Y��((��'�g�,�.<V�Mx`M�i�Ɛ%�A�D�P#���>v&�V]��K��$���vw�|g�lVї�CAtc)�ُƨD����ۏ���r��!������P���Q�l���T��"KXQTs`���@�e72�X����~ޠ�'"
\*X0��:IUaH�o��VA��9�5܀�r:ER�,8K��S`%�R�ϩ�n��Vw��q�o���%r8���q���+�ե�l�HAL4�����A�n+F�)iY,�ƥ�)"լ���v�0�*μ)���	�݆�m��W��(���j�Pf-Z<�#N�V��gh�{a��_C9�d�R�*N�І�B1 �g�%��o<���.�w���ʐ5�yǒo�Tn�# ���=�2��0��Y��=���Te�y��HPD58)���tv��c9+�3�쇽C���<��f�H0��Ȫ�|�I��Sc:w%8�5�e�RK����Ri*�DT@��jx�|&��9�@w*�H��d¬@B�{&6TL;&�Qos��8b��bo���:�m��s*H ��X A�&jd �i�\r�Y�Y ƴb��Xw9�y �����"�m��l�GZT��bv{�rKθA�Q.@Z�F
����-��-A�AYH�67�;�2Q/FNC����(��t!�RS����ڱ�M�M�	��6V��3IT��ȩ�9� �8iR�s I6�9�g��'�X��A���!H�p�݆��� D	=����@8((�U�z���g�t
�(,(�ƔJ�A`$5��{�Ժ=��/��y����r�M�H�k2_����m@/v-�������Hj�J�����p���*�`���+&��Ј��
ŀr�G�GH�챜�<��	'J��dX�]���g;j�^`���렒���}
������n5�]��#s���o7H�fI�ś���`�5;��O�l��~I��b�VT�R��?�@�B������z���g�/��0��@S|��G�C_ؑ����0�֛x�rD�
���,J��]����Tp����+=��%~���N��$F�B����!b���J�|�pCT8��i[쌻h5�-Й;٘�+*.��/���tpa��\���,�G�*u�*+z�&M��P���7��'5��a�C��*��A��B����QҚE��s%mN���AN�����W���cy�u "�!��a|���(�=�n�@�/�ۯ�V��C��o��x�ӍÀ0���8W��Q�W�	a+��R��*҃=f@ cX�+�l���c+������E���>c|?�9�L��f��{�h��2��a_!}�%�V!��8�*i����^����L�|y�UǇ8��Ė��b=�J�]\������Ebr�8�,K�PiM!��1�a��r����Լ��܅��Pm c�ͱ��^k��`I7��V�5�~�ƍ��׻t$��%���R�
�9Xc�R�r����hTĐ�	�p�?$��Ef\B�^�=��q8f��Հ��0���!�t=��7�c|�Gx���id�s$�I�5�ϣ�cY����D�*��(Ha������km���ё�%�-`�N�p4}�!�	� �)(���b��Je0��GA@�I�k��g�E�Ǉ2c����:te�����q��a�<r6Ո�^��b����4m�H�!c¤�U��xz����1������7{�P�}�j��1MB	0���K+����`P�#[���� S+[k����y�MP��{u«E��r�Ӑ��܃*T��`�a��f������1Ƞ���� ��Vb鈽#&(��f��b?K��Mq��`����<�}��D9 ����0�_ 
\�ݵ�Wo\`	
�ؼ\\�
{D�YO�'� 6OE����/��$�iܠ<�g��&�ZK�������8CVa-�\�x5��-{�����ǋu�U��3#c	��4c����K0Ҟ��)�tG!܋$�39��ԓn�I���TTt6��y"�q��6�J.L�ΐo���h��b���B�*D������kvMq�C�X�0y:��`���-��� ��xq�c;�|���}��\Yu�I�(ߖI>�w��o]lJ8���݃��qQ]�"�MQ
��-�bA�B������woOp�BN z̬�]^��L�^���$����9H�8��@���+t����AvZ�T9V�yz`D�޽{��ÝJo��\�l�Ve�b�� �(���$�7�Ҁ��_�7�9���pt0�2$��\���bp+�ߙ�P���E��)�Bu�%�:  �IDAT8���d����5�c� o�t	�ܢ�\M���+o�%�ظ��A���DӲ�������qؽ7�Z�5�Y�h@��)�^;�٥�S��2@j�Q�ȗ���<VF��Y����������SΘ<�䆟
=��မ6�,^U��2���r�c��"��s���+'��+磐
|�n޼�/U�R�a��� *�.|�s�j�s3�HĤ~���8�/���B�[X� �us��|����t�~��=dE*�P���'W�w�+�����oh$d�g��
�h��kC���0XE��>� ~a�Xi��H��qM�_�9�l������g���ˇ��$��I�0��d"7�/z�t����L��͌K� &E��[`}���_~%O'|݀��KC,�(���{Z��
*pp�9��s�
���}��W��o��Ò�N�{
<p ���d��ˊ��b���Y�!^��h��ǿ�^�J��=�hpm�-M�a���A�&oA��"OF���#)�Y�(�����̍3���tN>��lXLU�&�G~0%�6�U �
f�Ѝ;�a�P��.�;_���Np�� s����R����k,��~��|M+�ޘ�ʠX�k���xջ�����Koh!�!��a�ᆆ�]���?�����Vs��m�Z�J-f[U��,f>k
�L���\q`_k}�+��?��C"*����7���spTq�K��zS��l2�j�S��Ѩ}yRn�,c�	2b%�-L< ,H!V���?���1��{y+N�d���V�b�%��N��jjz���!�)ôl�d��'Kc!��;������?�;߯T봁�=ب�k���)��?��0_8@�P�֚�jw ')Fŉ^E��/�JC�S��!b�hRC���6����m>zP#�1N��)����A9�Z��n�67���#�i#�Pfh�r��V6$A�v��9���Q����F�Uk��~�Po�Zʞ�}�B Q �Z(�8;v��L�{5�-�XU$��䌞� ԡ��]�f�/N:Lq�:l�	��!�`��]�H�	ykW�H��
�+��3=�3����n�
p���M-�*��T�J�t ڜa���}� ��ᰆq�p�N�������6��b@h�!�=n$��o��Ѓz�6��B��$i�܇��s�'<Zm'd8��w��;;;$Ppwq���'�C�9`W� *�a㱗+���Ň�2�|A�u�l&
zC/�a�k�z��MR' BI�_�I��2!��a��V��U��9Q{ң�F�A9�F���f"5P�'0"��c��!\"XCD>��KɅ�	���(r��⠘�w�6.Z���AJ��_�`���N�^G�,�V��Q�U�e^����GbflE����
2�*�*�Y�C�S4|�K�Ds6kǪ���tTΰ�O�Mos���h�݋j�m l�&�Q}N�D8I&!̍��YbX!b��J���D��wC!;p ����d45�RB�mbl|�H�&!�'�L��< _�PL�}�xy>X$������KߤX�E���,��B�*�f	 ��$
YX���!*�:��O_��cD�Q��4"p����F�_F��������}gF��v>�
��$�y~y�$�In����R�g�677!���fkt`( ȁ	"�Vl*�= *�y+G�Ib*��8�pTb�����бJ�<N��Qǩ �Ȅ��9��v���I��5��a��ZE�fƹ<��5�z��k�?��Np�V�B�2>]�q���D���,��\�!�f%��"Nf(�s�� ��l�d/|��$�Y�������My��Q���I�h�M�s���g� �����f�QS��kKUR!��(0���!�a��MF���@���"����8h�w���7Zۗ�A��U|?�\��D�a�~����jg1�?}MI�X�hI)���ﭫ7c�V�j�P@'��L�b4�W���yũr\�L���Wñ=Īq�>}��3'_L��U�k��X�s�4�Y�}�H���PDkaߵפ�ۥ7Y��ԂKK�%� &��/bS� t����Ya�IX�!�ņ����u���`K��Cr�z55q����V�懟����a���C�,�p&��k�T�\��r]L�����Z}�]�%o��@#�V�F)]s�3}�4C8~���1���k��}�b���D�,��]l]�nf�FUR�(�W�;���5�kW����=g6@Z`���{��i8���pS�s���� ��5�f-lH^`C��*P��moo���7�v+��]�h���������.��_���#t�D����~�q�U>��/����y��"�J��lN���f�2��B�4V�tLgq�� �[#��i6�~�ri��~��X:h2.paT����_��0�=��*"�{ҝD�d` �1B7*�.�%h�JgD�ko�[��K�*U�=�'��{�w_��ԀL9LFxq��>�b�#i�g}CJ�l�v^�u:��^�����Z-��T�6[w*��z�8�s�G�?�{?�y�|���P�����C;���w��G_��ڥK{�]�D,lç��}v��t�p�i�H��4�Sfu1�G��e�C���'Հo�i���`��(6�����o^A����*Z��)dXĠ\FB���3&�*4*=���p����<�m��K�Q���4J0b<r���n/�z��a�լ�tHB
x�/�j}��r&7�8��[2�%>�#!�������͵�Zv�K	 �Y_k�x�� �:���;v�H����{�w�w�~g9����'��]�ɛq�i����X�{G
٬8�a�ï�X������k@�0l4{��7���j�U��7��r{G���/6&� ��Pt�+�1�֙�r��nu�}�J����V��'�j�mz��ԙ7\f��� c�s)G�:��<�'rN
��oy��t;ZRK�&���tm�D�(���`�YDL-S�A��\�0Z҂CF�Y�����v`؛zD��|?jOvV�_��i�[����[
��>}����(�����eZ�@oh���r�tз�fO$���LQ���Q=��M���b��uw��@�ڀ�c�����*O��ɇ�3�T��T<<��r����sM�o\��L^Y"��$���F��Ӥ%)��Ɗ�[��L����)�W�p�˛���݈$�uP��X	j�Q�6��F�ȧ����U�m���A�t����F ��^=�= ��(G������C�� �������k���z�r�g��9O�Õ���H{;���_)zX���8����ɽ�L5Y3ڙ�M�I���)Z�
 ��gkG��ܭC!�t�����P���d&��1��X{�#�N#�3xSW����~,�1���Z��{���<a�5tѸZ߭姟�㵝ӧ׀���Ū�\|���d:����ߴÊ�c� ��\�.r�%��1�9�Im��7����B�i�K�3�sK����֒6�K"��>$]Œ'$������W�=^v�l�lЏ�\꫖X�@�C�r9���y��]�G����R�^ڵ$gҥ���'}9��H�N���|�p5��d�h��E������P/E��Ա<�j����,+˦3�x���I��f ��<�߶������x�"�[    IEND�B`�PK   ��W��S(^w  �y  /   images/2e36d9e2-369a-4515-94d0-1575017f862e.pngT�ctd]�Z���muԱ�tlwl۶:�Qq:�m�v��Kw���1�G���^�=ךs������8�   ARBD  � @�AC~]�������p ��}A�x�K�.�8*��&�N�~��
� 5�po� ��������E��֑��k �#�:�}��E��h�5u��T89�9��}1�y{�I��|�7w���ݱ�,��IG-n��z��yk����}�|5�HrE�;45�uA�u�m�Kq�^ ^8�?�����o�+����O5q��ia�tv��I�V�qI���` ����79:�ٸ{^��V�Y���\�~�}9����S�U�m¬��K�Q!"���g��zA ��c��!��M�~��ٔ;+��f�M�'����;� ���	�$!�x{��&��.����݅�`�M�mQVN�B:g�޻K1z|L#_2"1����o4pO����n8F��D�b]/�7��i?�8���9z�R��H8��TjU�y�������+�U�W|t�"rr��(a�K�w
d ok��{O��.Q翤l#�5Y������O������!�*����r�AE�����!���Q��*+RQ�Q%���Q����}�\�T4�\B!�@^#|�pAʉw_���<�}F%�ؑx�\�����+\7����пAQZ>"´?����@h��E�)���c�&������͒i�2���/�>��ɺ��]�l()�bt)�;(NyE�x�I&J��\�_+E�P�;��^3�j��ώ��������_I��/*���߀��J�����0�B�ɘRd	:՚tхs��Z�<nO�]f�[���Xۙ�~?N�:�O��2tm�ݗ��tS�6$Ҡ��d=��_��y>��>��>��'�'K�B��:i򷮣�s�[���c[D�8���IK�3m���$�5�Y�:�E����_�^�!��7�<<Q׫��Ўձu��Ixڪ��]o,Ss�(�L|붨i��X)t�mC�y�B���T.�D-��9u���2i ��n�������x;��T痑k����R����rTA�WZGilO���\j�����p���=�Z�
��A:L/;��m�,�h���D=T�+�9ګ��[�1��.SRRJ�YҀ�^�-�({g�J�D$�r�����9��ξX����?g�d.39�L�:��#�"�I�_�d��x�@��\�b�L]�z�����������w�srZT�t���V��
��t�P/���e����,�P�J��5	O&�u������&<i�:w��:W�O�V�������t��ݵ��Q��q���^�YD.�$f�[R0�v�Q�*u�Q~�/둪��LIP��޻�� g�8�����bw��
�K}K�W���166���@���z���/3��&�K��	cz�q'C8��4����s��m,3Q�� y��\*����){�999�%���<�Ml�"�t�z}�Z�_�5���]c�����yld$ͮ(ۑ�kc�))EWM5���sJ	���7^�����Һ�OfG���Vd�dq=��a�!,�8H���� ��P�^��-�\Y������)&�n�!�����I��
�������Ԧ�����@� �>�}�Y�}���)u�k�~�B@�[~!�#�|�)�h��Ep���g�	AA�NF��nv�0 #/"�?e�?�#�hYm��v�{��k9�n<6aw��<Q��߳U�fD`4�A�s�>.����f���5ө���C��D,�z���s�:.򱺼��ש5d�*«l�AA��s_F�F�$�ad��o��23�7Q�ս�ٟ�=�	�M���\����'�׃�^^���}����?�39sm|��Ǧ���];=�Q���^�����k��qȸ��Y�K��Um~���,�z�n�������H<��_���ה3i��m=����������執_H!E����;�]�e��w3� �q"��ADF,���������i��<�Z3�f���V�PY���ӂ7�٭��@�S�;�d]������m��[�0���/t��V#����zf�0]���U��r�q��1Ja�����
^�|���;�*�W�*PLvV�Y�0v���|�����1UUҭ�ݵ¹�.��Qg�R.�^_�Nig���f9��ݜ�]�5B����~��4��Vg���W�IB���M�]@�B���[YW?ƏgBVM4T]��_Gã��t�2,��1�WL�a�Y/O{��2�{�����1�8���ʽ���J�#-�R��%���'����-=����{�hJ���Y�ݹoS��Nu����l���GޏN�Ó���X���N_������CR#M�������f���Q�h��:�q4,�jT���)q̛�Y$P��Ւ6����܂	%���zt�:���w��R���?����/��B9�jʦ������F����P���=�d�e����L��v��0��.�5�ӕ� �3��YH��L�}{xП�#�P"{42�gM�9�d�OX�3灢�G�+�F��H�dv�+�?@�]X��=o�Jh�3�'/bJ�Cߧ�;*�*4��$$�M�y��nk�� 9�f^�r4�;|l/5�|���r�
�x��`�2{���}���JWFA�=��+�~�UT��'(,;Մ�U�����ES�-=u(�\ �Il�Ҋ.����~ǣO�����cǑS��ka����G�r��NLp������@Q����KHOf�٫��+��@~.��?E�<�l9Lr~J�-DJ����!��g���k]%ʳ���A��{}��v�AZ�	,���!Ml$�4�kބ|���i*�rk���`�q�J̱ȼ������~�5%�� 8����M���o���.��l�ח�����e���~���:���n��|��[0��Fy��{� ν�8�VR�7%�>D[[���P�o몐��A{(��;��:]UOكXE#��I��נk���)6����5�����;A$n�3aKlL�>�HU|^q��O>U˽�V�x��d����᥆r�a_W&3C��<�!�T�wJ�0��_�ɛ��#]y�Ԃ��y~��r�1�9{z�72�K^�l�W#� 6�^�9ɖ�N%c���׵�(u����ZɏZ}��f	v��KWQ����+.��f �!�w���f7�>!ۇЫ�����唤�+`���^4m����l|�K�x��u�D�Qۏ�,'��s��w}���I���Z#���v:�+;�l�^m�h=x��M�cG9MgZ}8̳ ��9�r
��	W���অ��k22;�]��,8�/�;����-��͗�L�rR~�lk�0Z�J�����B7v�u��=��>��ð�k���N9N���g\���4S�눻Ҵ���o��"���(Go�_���V����1�f��^VJ
v�>ͳX.\�W�+tN #!�Szr���sAV�mĭ��`��QV���O���v6�A%���1^0�]�m��j��)��=����pq��Q��"y�%�NG���X� �՟pU��9ڱ��+!%��������'����BZ6Q����e�#���hf�)�ꂬ2!.NR�����`�iI:����L<��å�"��\V���5p�<s���
�ዴ�=�޹&s$�i��![M�K���<�\�n�dH������<lAR~��b�7lG iI��ZQ�O4B��ƿݦ�
���ءYվG������b~�F&
�#b�l�u&8a�77��S����,ӮY\պ�b~C9p�!�a���'�!�$e�w����O���Յ�����x
s�Ga��a��17O��+�d;�+�G�3�S�U����+֟EWO��J�8�l���� rG��D�l ���<�4Su�at�d��ƅ�	�S¬�Wp� ��2��1k{+���PfNځ'�At���<_�S���fR�i�, x�ɯ<�����Jc��H�3Fx8�l�*9�NV����&}�`�������Z�.p�z
�Ωaț�y�|�p��������JvO�P�3^�<5Ɔٻ���o��||b4'�I������~�s)�ښ(!O�XD��JS�^V��7//V��ݹ0��(���������J�3-��eUI�T��LL���ll2\]�lᇇ����(�ӪW��F���W���a~�4;@$j��*�T����B�x�$���+�g��?'I�rb���D=��,�ˋ�ʺ������n&]ي��x�[� �5V`����[�ꝕ����m��$;""������6�)�_�uH a��Hkn��߱;O8\O���c�20�((������)k�@!oJ��lyŞݟ�fVX��ך�~g	����t��t\VC����Mz<�~zeEE�16L ��ӟ�q �����;����Ѝ���q���~����.�݊������[<��"�8��Iy�oJ?V�z/��$���݋��.�j���XZZZ�������A$�]ώ��^g��+�5Mun��uyy��a��6:���i�����$�w��+)���b>×ϻ�����Q�^�<�	G�c1�����0�P���o �Uw���*hIs����ott(��!��Aml�q���o-	k�ZC?����}$��X����������K$[UN6v_IL<^q�w�O�p��q�4�"��A_��š�4ť�Q�7_�3�g�yt�z.=\0��=ϩZ�-�,M�#5�w>�y���N�){O����L-����om��-T+e#��j���@l�q�]�'��f���z��ן(��}PQ�����@�,�^ػ�*�l˼���SD��̝��ɰ �RR�zb�/�W�����=$��#o��hP�'#��ğQ�ha6R�Ro���l�:>]}n3���Ay<S�f]�"��1��� 8����IԔ�B���٫/�@l�'�j5��Hl�9��X��ߣF7<�|0�q�T�j�� ��&�����b�X���BQz
d;l��wx鈳�pZfz���\��&7�����F�k
:�Z�#�t�_�n,)F5�_�z�O|;A��;�s��g蕬�-j�r�c+�r����>���FKssS,EH���Yc��:�z�j�_w���`����^sp2���͖pP
�ֶӥ����Cp0��~���Q��� �^�M��	���7�3� �����_����=o���ߏ�v� �!�:/�渮�z�X��5'Hk�~��@-���^��o�xM��'2=�ЗG�o�,0�i��!(NZ�^fO�-Ъ�-r@����4�OH�ٓÙc��8E:��H�$���Pѭ����Ǧ|^�?Wk���ܣYx<���ȋdq1J��8��y����~8<]a�po��5:��!h
�*��@j������j�*��֬�|f怜��D@5�*��Q��Gv��v~�&qz�V.��߹��$Q�2��D�i���}�>��,1�4W��>4�q G��Y��Џq�{���X�������I�_Wߣǒ�?��*(��?��7��X�Tg��p�~�VZ�ƍ�O�#v{���,%�8=�WX ��C�C;�s�����R5㈬G��?��{�N1;
���fn��x<p���X�xk��z�Ͽ��S������}_M��.�p@˲��-&^	�������,?��p���W����`��C��s s��M�>�	g�7tI?�//�R<2��`s�/w�u)��x:�2&f����;.�X���+jKf%J������M��6���d$���.n�G^�]`q�T�~qv�]%�ڥ�UY�U��acX�{�%{��[	7?��D�	���f�Z�?ӧc9��D�=�	�`k���Ͻ�H69g��J��Z�#��ȋ pr&�u����Ӊ6�;(�"# ��5���֜��ge$\��/�P�:�s��3_�c���)�>u�v����Q��+`���,$���X��0v��V�i��X�IwF�_�ši?��l��"A8�pu�s�=l��$��l����8x*��y��٩�a�^V��Ho�эML�>�s�XD�XY[W��N�"w5��L�7ʒ��bZq 
��`N��n%�M0Pz65�58L>��Ҽ:jq�Ο�u��  �b�\��k�ii���Z��l?��u&��~Ϡ�W8���,4(��h��j\qhjBz� �@@0�g�м� !WZ��K�"i�;9�:gf=3*X;�a`aJ���}b>u��9s�e>n�m���B4�JA�o.~)"l�zlS
㱣L�^�b�����벛)�1ؘ[�Nv���uP&`�S������.;6Ek"t�Gս<��pNɭ�k�gEݾP:?�Iݗ�c���x��	4������Ƶ�_N���3z�]��]A���籙<R��Լ&s�����̙AR���f�>� W'>a}�\�JS5�|�\[.!%�1C��z�vy2)+k�1k):2��ϑ���y����c�P]�Ɩ}�Nv����c4p椂�m�A8rK��z��+¢�[��d�!Cb'9�����tB�h9ؙ��6��nO�[�m�d��mp�Sg�&/�����d2s߅R}5�'��l�</r���Y�Q���vq&L,�
��^�>O����X�b��本�\�����!����]��Gܚ����̀��� !r��$����{��}ۅ���n���B�š���l����27�t#�W��J[k�q�.�v�E@67��e{;�$�x�E%���M���ސ57���X�|Z`���U��u;���ڦVk)9�9uT��"����ѡ��nY�}e��6�Z�K�T��/{��v���=�{��pkbJ��U:i��[#+<D����B����X
�)*^�9s�5D�/}�Sd�X�������|6���M���E�i�=9��S�!+x��VT��w�7#�[��͞2�_֝[a�	��(�x�����p�925l@U4�+�'��彷e ��%��V�렚u��B����.���U��&B�,�w���wVJ�Y��t�lM���8���[ 	��@���*<�aC|�|��|�L�j9pQSW�Q���0x?��ፍ঺��Mw��k;����/�qC����/oa:5s���7�������ra�A ��ec�*ɯ7߸�zkG�L���ʳ�� -�sVs����;�-.��H>�CCC��wT!{vg���9�bt�eXQ�����5��9��@#���B(Y��)��Dq��ܡ�li��~{G,�C
��������.ij����֫�Ɍ﷾��oo^��볞?Et��ޫ ��f
�eê1S֝����97�l�L�t\X�@ʃq�=������_;$6�:vfk�g�asC1�b�?�6��7��t�����IY�X���*��:���JB9�nn]��4c���;
x�
y����<v6p5��ҙ�v��w���+���5���V,�����GG�����#3�̛������'ݞ��8���~χ�� ͹���Em�5tҭ��H���Y�T��r��Ҷ�����{'+y����M7��ʹ��X)��Pj���fN�\.~Q�rvN������
y��(���ޮ�� �k�I�9�ϏOG�&kq|�\Q�ȞEP�~�,0=(9�:$;�6��{���;�g7�~�i�I׎.=��q�?������x0?䆆๹��V���=/���_}>�P��Gw1'T@�����&��B�[^��fd2�����pS� }���.�,>�֊��vp�q5����IkP��uc�qsP$�F���E�-��%}9�Q��t�Io�-�p���KU-֖m25��@�+x��kv�~H��D���+/�{.aj��N�BK�	���`V����1�^-��-l��;ޯ�z�ա�r���g�uf u��W�Z�F&�(���%��DE��h��S���o�β8ֱ֩�)�s��Ifk���+��߫!���-䉥}����.�n�A{p�!on^����M4�V��(�bK11>>��`@!xcst�9�,������;�]� ?�$�v��XRZZ����Uٶ�$mH*�g��N{����o�熹���~N�[g�}�v�h:\������-U�5��̘f6^_F�����C��)�GF�N��rf��rr�K��6J�縗5�26
i��WMpc2�m�+Q0��nj:ufk��ݲb��ܔ�^�v�,�ߌ�͓���]��>��Z�K��sT�f�5]�jg��5�N�i��Z��%��'݈�n�7[�}Z��`����n*0�clFp��r�|l���ʕi��T�[K1��5蹇�';K(-k�v��w
�';����GG�,�ҸMܭYwis_2|��l'��H������t����71?���޸fT�QP�պ���~���%����0���W�V/vd`PejwЗ0dl݇��+�+^��� ;Fî0��/���渁y��H`wK�5�#�o�=p�"�&&�t�K�Pl5�9��Q|�$+A�nw���y>,��<P�@���$���K�M(�GoiA��
&�UX�孪yW���"|�C�<�5@��J�!���*o����N��?`�	\fH�X��{C"A)���Y8��t���o+��xj+8N����A&)�;�����i`���۹��p�C��:����DbF��)�Q��PY�I �Pf��R����4�(mIq~��(��v&]hhT��+~&\��B��a9նT��eIb@��K�CE9����}CH�x7.dA����'�m����x2�[��7	(�'�G�a�_9]��������R��G�N����]m��Qe�&D!WTs=|1OmhSD��;wV��nT�ȹR�?�#�����P5��b��7O������A �p�w���m��k�+7�%i�!��u要��L,ŭ�@w���Ɵ+{b��L�O�w��d�o��5N��r�h�22laų�a�\r������k���^)#֯���I��S��=����Y$����#M�Δ�������Aƕr����CR�z����kV���1���ڐ{���9�U"�kOF�$�������]�mgn�"�������X�7���n�E���d[\XHHH3+/��wB���C|ߧ�-�	#z-��o��ѩĄ�ڝw��h��`�m��w��+{�ޖA�j8y��\ݧ'>�ˤ�?��[	A�)TB��L14�i2�������xP]��B�$�p�I7x�%�W46�+���T�%Ћ��}�����(�'�)2�&J)2`�{>3��V~_�
�![�(����,�I��u��މ��3'd>�~$���꽟��/b6�v݆���_Ĵ=��1	��ә(���)c@�u���K;�8b�`��s��O|��!?T�6	e{�����t�8�?֡%���FyH�X�j����=ujt�ՃnJ��n��r�a�9�LxK�p�OM8��K"X���#ˢ����?mjP�x��7��j]���/��}���8��� ��޽��T�����dt��شờ�K���)�u?n�~N�v���m�ǋ���ɑ����r��W"��v� ś��h"�j����ʔ˭�6ev���-���M��� �îź2�5*��Qx��֝�#�,��Y�5d�Έhh`�5�R"��K�/�Q�?>�YߞĞ(;:�Ъ�~�K��Ε�錧��7픸�k��/��@��E>ePm�SL���'r22d�5���*�� Wf��R�����/���L 7��xH�2U��
�}�g$ r6��6`��7�뉧�k-�YQ�U���h���X�[m��B��qS��3�_��G5�஭e��ZXX�����8x��6�QV�s�a	t�m��$&@��k]�D�����y~G{� ~i&��/���b~�����ť9a9�k�$5eŭm"��(�16����-�C9*L}��B2^zzz%";p<����_ʾQs��u�^��|�b����kV�^fU/M���y��eTP�@T.;F--���g{4a�y5%]/�}��? jsf��˥�-�;�s��s������xk��&?�w����M,�@�v��	�P�*�D1�3u@��?�H:bm�Z;�g�v�H-ek}9�N�M���!�����`%I�L����&�Gpq��k�0�'�¢�,%̔d#�0sŷ6�FCe	FFzT@�t��>�(qVn�;���PBb�DޯˎW���{b���.��;�8$�fj�U͂�fu�~#����`#���6�BaXvBf�8����A

h$�����N�b7����-�&C���&��R}jW:oTP�nv��B#0|��Ht���X� �/��>6�9O�X�^7���)��2 #Bx��+#����a|{�{O��i�����( a��ƖTVV?�O/_���_��X �bx�r����C<ܚ����\-u
��(�AB��􏸂q%�.�?��pT��bu�<?w��It��Lc�Jw�Ad
#�M��)/G �2����J��k���5nK0��$�)V�����S��ܷ�#3\��y�v�g�C�#����ʯ�VW�c�رa��ʂ��G���C�J+D<�u����[쌝�2)(��N�"a��j��B2%1���A�v��i٩)͡,&0�m�Tx,��3�˶��݇���ݷ��NX/�n?�ؾ�0��u��@�l���>������ nV�nNY
��
v���0(�����R��@��Y��V5��I�]�O�)g}�z�0:�:�£��w,��͵>?w;���eB���g�d�����D58�l�NN��킕9S�q��4��+�-"B��O���Ryw@��Yl���5�\�Ԑ/���1������ɒ�` SO��,,�.4E���1�k�?���O'2��f�uΎs7;}VU��SC�Ғ�`���Oi#K[�`�`�.�7�r�춎��(�0�,X�Ӭ`�����R@W����1e$������D�r�c�Ծ�b�����ܱ�ňeKG�$��Y�:8��j��R@ٕ����������䚸`��q@ѴM|�����=��:l�is���M�D��a��G38�i���o�7�3Q�^����/w�7���%U�!�[���lr�U��t�ύ�  B{6���yb��9J��\�i�p�1���h�䉝ŰX".3�''΅���I|��F$0�k_��[ܘK2y�Y�`ss�5��˭�ފ$�t�<~ԅ:��S.�nr��o*ތ.f@V�D��2]���I��8��sd|6[}x|��=I~���挱�K����bO�ϑ�	s+�� $��\T��{�@J�v��i�,��=�P����]�I�����~# �I2Y�Ҋ�{p�y�y��s��e  j��]��q�E���p�h~��3�Qc��ʶ�������f�q��=�>ƒh��'��^�@���Vk��D�-�܎i�7�e.��O�m1����=�����������(:8f?��r�@��H�y>e�>�C�@RBJ3))r�������Wr¹Dh�*�0Z�l������RcD\�c�����;��$��L�J8������֏��2�܅�&���UTTD]�'���n������m���jk}�I�R<t
y�-�`ˊ��jLI]�����0�Y�h~�RqL�E�a%�~N���aac�p��fL���9f}�KʵNgp����$�)������m�]3����w䥁�kĚ����Ξ�����߭o[������G����Ƙq����0���INFR�|Yc�щWtK�&>'I������;�x�X�U\.��v��_m^l���وT�:�t�1��SD�0�����	a���W�ц��n�=(�������EKOU+yO�ϑ%��d]�!B�����;0�-�`{cɓJ�OsH7$�OCI���\��h���d���f�~���u	"b��9�� ��<T�5�0BN�%���M��#io�"�f#5޼�]!�
 �S�f.�ϽT��1�;G�c�W��#G&qS���d�` ���C� Q|��r�Me*�_��j�tM��	�fd1\�z�Gw<����r
��6rq���4ƕUTQ������."GF�c��6�#zqNj�i_�Y�	�o�<�K��޲���?	W#y�[w�P�!t�,�#6�,G\������]��\�<�&����^+��&T�'X:�ХG�C*g�Mr��v^�ye���A�.ɕ%`ܸ�"=��������j��U�y��bx�l�h΀u���)}��Br��P�~H0aae}�I�m�L���i���u0��c��U�s�H8�S�'��K�A�����yA�����r��I�T�¤��Y�����Z��w����{ ���c��D����R�2�m."rNK�18^	0�b�<d�Y{譭����P���RO������mb������g}���ř9��hU��=m��F+���Y�
B����_a�@!v����o�z��-�'k񟠽ͩgʹ?���@7�z8�F�=��w8����z�W���dC|||I}�df|�M�lNZVQ�����N�A�|� S̐�Cٶ!��-u�����U}��w�������ff������X��M�����'u��V�!ϨG/f�M/[#�حZ��M7�)�	��;2���b���d�,�?�4��n]���Z�Amd���6Z�	�	Y�Ͻ�v|΄2W���]F�))I?��i}���X1��׳!��B��+��=��� �����~E,�����F>D�ˉ�V�E�Ą�a�{xV�p88٨�ar��$
ͽ"�vX;Y���1�iG�^��F9W�2�79���3nFn��Pj�o�_�aa��.+k��o�ϺF~�?ې��l����YK���/gm��p��5Yn4P/��ӳS�o�ǻ	ɪ4�4������թ�i�nAp:����[�Zb<BB`��b&@$=*
^J��fD4u%M#bmYm��q�e�͸b>;�=,�'�ߗ�Q��Æ��_�����^ݗ�EUi�-��5Ϫg�]b,,&����&�U����m[ժwo�^�oZG]��������ރ�M�/n�JI��h
u:J#�y��r5sK�8��&����xE���QF��y����ksֲ�&y�g2\4�y������!�W�^+��݋ �������Fv�G_�jc���a�.?c0��*�#���,&gU@E*�]����e��gS�i���x�E������5���|�Q���}'�q���T��6)*ʜ��Q����!�M����я {������$��>Φ`D���k�k���9=Ci]���+���ʯ�1�6�%�2����߷MZ��L:���5���d��ښ��~�L(=���|�D�i�Q�Ea�	�C���|�$�T'S�w���0��D<&>��A�1��� �p��M�oi����et���ղo��,�]N��u�}3};&<1٥��uw��9N�Ь�RU����!?/O{�T�NN��}*�\__�á�Εu�ܯ�*I���x�b�2a���ŝ��e.`ez�#�,TTd�Hԉ~��u���4���3����Pϕ
{��TN�i�i���9�[�ԩ������cBU��-j���[���ʝ��MK�2�v۫`�@���Vc;��`�)%#�%� �`X�5��U����N/N,�	uk���wE�J�az6���v��V&1�5͋)� HI�i���v�����ߑ����A*��4��r�ڳE��3S#�����Dy?,"�o\��Ն�8WV�<j��Ayz�&��</�Vn�yW<�|�G�9���2��kR��K���#&*��B|��nr���;��܉ Z��:� ����}iiIJ�]7��t�N+f�Wtƀ�x����cN½y&���ֳ2軦+;=]E�۰���*=[��R�AN��}�Ύ���s9��{�;��\�I�_�$M�o2��$�����-���'�ɱ�C��&�/w�n�.���*��v0]�feDb� ����קI����z�A���W;u�^���]���FH����_W�1����ƀ���^<<?�(�_RA���]/t��2���[/�ҡU�,#���RQ'��Z*m��kt��Y�	�A&�ֳ����~4������3J`�1J���l++-�8S�}�j�,O��� 1���?�jk�Tò��\��Sw�PF��V%(M�)���! Ȉ/�!��Cd$j��dab�JDʢ������`A���"�t�+�.�֕�¾I)�u����]�Y�d���(( ��!",�ȽZ���3��d�wLp��,��i'��������M��^�\��
�υ5n_J�2^S��v�+���
M�3��L���j"��ǹ�!���V�O��2p�D�Ӓ��:T��n3�gʜ��C�:&��`El�(S#�i� �_��8�%��h*�m}x���l���*��i�hU����r����%=湏})�lE���Mۙ�=u�R����2��#Lw��RR��V5�o�~_X����Q�U���d �P�B|�'n���ѝ�Q 3�X�72$s���DŅdcʓh�����\o��'L�6R����F�q�q�snK�X�/R`���.m�����/r������ڄ�-��I��|�rÄ��~}XM5%�S>-��3�k��N�   Z���A���N� �f���o�f���m�ҏ4E�쫨���!��L�s�����r�^Q!p�o�ʶ�W��iK��h��:�v�3���'�v�2RZכo`��>(�6{J;�S  tcJses�����u�@s^Ig��^p�B�����ٺZ���4U�IWEm�����<�?��9$2���?�������ͳ�g�'-������U��o�E'^�Zv���'܇��:_Sa�J��j��?��D�p5n�K���:񑴞��,����ǳ��L�M�Q�����cGW����!IWw������P�<lV)��dk����G��RBP�PSlJ���P���}x�e`S7�TB��	��3����,�{Psrڡde���|I��J9��6�%h]~��AL��t�����~�Ä�ciQ���v�J����WYI�dH(I�_��n�[7O35%��ԥ����ͺ�����=�RC��\jW�h\����Qd��P�1�w
*Ε�~p�n8n^g�gػ����%p���A�� �����>[e-1�9����a:oBGN��:���W��#9�:���G���۟J!��S%����Ұyy����̗��N��mѺ�8��B^~���R�hQfy����\i۶�P0��+R���Bf���/���˛?pW،(�iάS��S�g[�b��E�������� ����r���#�=��Z��[ A���j�q|���H�Ģ-��s0��$��`��G��}�ooP�3�5KR�)�����S��n���i�r��7^T�`������K
5���+% ?E���h8;���8�ha�C)��13��rDƷ��e��]�gL�o�7�ݜ���M)^��n)��!�u���WjQ�1�����3���]��S��!��h�r_W��85�0����o;(����;#�c���	媧dd�tҧ�Pú�� ���z���Fľ�ҋ�ۀ$	3���wͷ6K�UN�=B�/�n�&��{�NM��B���g_�uu 
*�x��R*%�Gc��
Ju��$t�����fF���g�I�mKk��G����S��T/�����i֐W��V�.^|���hw�b>s#ٓG����쏖�3��XE�����Q~L��+F��vA0�3�F�2m��YX�X�����H���0n��(8yl���m��(��@3I{3�j,_]�Y=�*ُg0[��®�<��k�XXf^��pH�W�7_�����\{_Ԯ�|�\������<������%��<���MyV�YY�/Q����5b�?(���Ue �x��l��N�QV�2A��4�պUЉ�	;}��qmZ�����<�d��PggEٖe�1[���o�ـ�!�ޓ��0�U������v©5�9h���$i��@��g.عD�X����C�Q8U���n
:P�  �C���.�毤��|k��B:W-z�!���<#��JVvw��]�RBz~�jv��?D���J3:JMI9��>�Ba?�W�L�aN}�'F�$�SC��z�)�	Dб=���{� 
�N]H�;�t&Mn�j�F�+CÀ�+�(R�I����������zL^������v4f�o	���h1av/d��=N�B��Sa����|�� K�?!{?�~�y�[���u��ϗȜ�񨕏v	px����gN|��=J9�Nb�7x,3G���	�,NWUL��9U�>s
k�Th~{n,f\���C�b\
h~/��&���0�eZ��RH) �J֏�KtH�z'�}��T���iϬ�@ؙ�����3X�E'܂[p��n�-��;w	.�%��@p'0����z!�����{��w�����뭪���WH_��^{��4����K��&��B9�吡�wP���vD��?� /�b�׽V�����Sr
�!mἓ嵢�?�?,ޭ~�͏M�><�n��c�q�Ko���V�>����)p�[��>:Iʙ���U�D<�tՏ�����+`-BB��4W�Y�MH�AܛM� 
U�
KGmt�mv�QY��,(�[���6gr���}���jR\^O��>�;0��9>?����ak��k�M12�4��2$��Xo���FffG9�ý�霞��~k^�kfN�1
����l���޽�݁"�V����I�G�<J�E�1��i���y�<7B�{\����(�;Q�!��=� �_� �:��������O>�y������,�0:	_��[ �A��Lsw+�.)���c!�E��x~�`C<]_7��JX�����^�Iԡ�C���O&-0\����E�*V��tE Ҕ � z��Id�23Sq]ȉ(%ɯT|��X�FOlc�n"��%đ׌5���N��'���J�<����aO1��pL���V���:v�N(��������jKp�؎����j#�%�7baa)X��d=���d[�����;+��M�$�c�313��D�׃��০ap��g�i0��OfR�$X�E�2g��Z�Ĵ���2H�v�F4�E�O�����	��q�/�g.�B����-o:�G¶�!YLzֺ���r����3Eyy��U�N[ߗќp7�8����j��͈P�/Q篸�Rz�	�jIt7cL��~����J��3�Ƭp����mb:q��/k������IqyY��nȼ:7`,6f�L>"��j�:�ڠ`fV�`Ғ��X���kA�U�bF�TB�xD�'���n��蛚W~cao^ _�x��Ɣ�?KL|R�ظ�wkx`�<aD^=|̽�<��&��x\)����c'z����G�g7恡3���bg�ȊN��ٜ��(�1`�����uR��2I'<��w]���lݙt���ż����Ȑ����Y��np���\ed�قM�)�ת�~�؋�`�b����e&��h���y�UZ;���m�:m�^�Ϲ��*��cէ�8� X�'��oKC�G&&U-S��5�����Ø&�M��&���Z�W�R������c~
�olI���(��������k��Z� �~vҰ����`�j�-�p�:v��5yvx^89g��6�|S����@d�R� o�l�碾��� r?؜k�8�&�9U�s7�y����<M����+�{Va C�5VC��r����`��ӹb] ଻8�&󃫛����	�1h4�Z댸ra`��!_9�=�h��$���IV$�7�!�6'�00s��X/;e�}̕~#���r)j��!����������e7(-���oݏ\�$��o�@-z�'$���2b���3owx'����t�P�n��J�Փh��44<l���xu��>��RDt������Q��x���jՎ ����5��3!�%��9R��Ԉ���ϫ���O@��$θ�W�6�%SS�X��͐QҰ�����p�-.�pf����y���{��4�z����FΙ[[lJ�K�.��J�!�p}�K�ͭ���'O3��G�Z֭w�Fy�Hrs��ib8��XG(�Þ��>r ������
��d�}L�
ځ�O�&]qVY	�4b�zY��A�����oE����c��u���ϑ�����r/�/���3�ɻp|8E��|S�w�O䁝���?�	�2	� ֩�ߚ��?�lc�8��]���ss�Y�f��9`jsߡMP�@KS�{s[,�+b���0�L/#F(������o�����{o�!.��\b�Y.�=C.�  �𺖈��._,Ҧ`fm�����[,����� �IL�]���\vr�i�ǯ򫪤ܺ]�CM�h�z��y�����=��9D"j��?׺��b��uc�@�vGq�M|MV��	�(,.�>vv?������>���G�|��L(�w Y��r���ぷC��t;rQ�i�C�ښ�2bE��������m��1�j��X^����`ׅgh���+<C�o�Y8�G�194�bKM�'�6���+z����.W=�v5^����OF�E( ����?s�ǥZ����[���nC$������ٕ�E9��B��T�a��s�/���Uu���}=U��4�R��&���z:�Q^
�T����=Y�J����7iƊ�vw���>�=V�"~>)�ڠ���xƝ��ۨxD&4W���n���� ����$�{�>_���,sw|_[[�a�"�#�@�<�aH<�?w��H4J���BUǛ��@'{T��99��,�s��������[�]{�x�@4^i0�}�'�aC�=�\������yNaz46���ڊ�M!~F@"�(�����+f+�Բ��o)��x������î�G5���.ƻI���3\�}/N��k=�m��-+���v�>��,�|� [�1���#�(�2��������-ϼ��@[S��R+t��x�A  l"���e��<��{��.��*����Fm�(B[���Mx$:��P�Ҥ6'.:]��m=ȋ0Mք�91��1srR�Xb�j�%��d�`��:և�ߜ��qxp诸�C��pg�`����c����H~t�{���̩��ƫأ�i/o��	�S��p�?{T���>�<u�Mϱo�B :���y�1�e�>����=��Ox�Zs�26B2y�y�����h�G�E	i����������DE�<C2b�=��������o?���N��:8��TU	�ǳU}������t, ��+ąSU�j+����`��#}݃a�)�<�g�-6�++��k�	e55,߫_(���q��^����L�&����+��J�BnZ��ﹿ�8Up�pA7V,J?��v��z�gFs޿ f��L�2
ޅm���G��`��#cUA]��Q���:�@mM��oA EW+��kk���ņ�ޚ<�;_(y��\O�,/�C�����"L�v,�s�}����<s� ���ۻ#� ������x��Me^�Ά��v ���`wO����(<wS]Oe*�h�`[$�ʙ�	�F;���`��t�t���5�)dd����yc�K�!��v�sҀ�����֩G��4z0��RV��C��m���
+A�(��+g�� ��$k�ߗ��7	^38�۲7�QZD�
�RRx���Z%��5h��V5S�]n�3o��t��	{w�z|��৛b����a����w8��w�21���`ɼ�e�͡ߘ� *{�:�߅/{��������Z�/���b�@�2�	?`��14l�Ќ.�T8iY�H�ȍ.����%)([Hd  /��J�m<{."~�(��Y�#~�m5*�~ ��Z�?l@��KQQ���������*���^;'�z@���e/�
�*e��2��K�FJ�*�˩{���h3��^��X�(�}QI�֍�����߄r�$������&���Q���}&t"sM����_��̇�p���h1�?<�Mk�6�T�'���
<��6�N�w?R_�����y׃�Ǡ��y����I�jy1��}�ǰr@��Fi�'���ۅ��Gȅfc*�¢a�!��?K�X{���:���5����r��%T4�K?mK��Pe%ŵz{O�}������λ�7E;R��s�)�<_�8c�_e~1��_��#�m@��{���''A�=��|��S�а�bU�vӔ�nD�4�į瓰i��L���\�[_�L0�/>�H&b{JK��������MA��H����^&&�y;u�o�Ϩky�W_u��|R��[m\q���?Y���=�� �sN�N�xO1��6:�+���etሼ�6���v6�A Tö��`_�3|����+(�$�GY֣n�p���NW=�ca�����}�P]�����:r�����m��O�����0!�a�*W@6�`}��F?��w0���^jjq3��Pp�Us� GJzZ���[|b�0$3_�}�T����~C�^Q)H(�:��� #��]B�����#���i��?�O�ۗ�#��;����1%���)���T+�f�.�A�������T�߯��$[@C��3X����k�A�闄��/�2��
�[6+|�X|�8�0�>��u����_0�&Z��P��	4Kt�ܡ��f,��N��10��d�LB��c��Eֿ���Z+]t�����)�/�
����tE����=�M��j���N3�L��t���FXZҼ�nEGW�gd$mZZV�]���s�df�����h*�E�9��zH�V�&-ӛ����!B��ly��Mb0��8%�V��z'� ���_�C{��˽�é��������w��0!:� �);�Xh�Aɽ�_���"��n3��بAjs�Y8��5���~`po�X���l�.�� ��{u$���2ī{�֟�:��zסh�Na]�Ѽg�>���>���ԗ]�d����"�q��T4�TaCô�Riu��W�/8������Ҵ���k�����4�0��hP�j��(�>�śP���}�sU��-�,��Jn02��t��x����qV*�����{������G����
�͙�I���:�D��#C	�W�o�������g����������{'.h����E��x�O;�G�p����,����q��~�dA7�}͕����5�n���a�82>��~��� �s�3B�ӕ�� ���08�,&b��7��ꌣ�e�O|bx���5����E捀0.qz(Vu��M�_޿����C�n�L뻓
�$O��,�%��o*��ż�-�:������|����i_���u�B�O���S��3]��$��xJ*;���1�����f�˙��|��Q��	Sp,��yKkkqw����U圞�M-FN����$ARŘ�����Mō	!��Y�#�u�(`��67�6�ȼnQ'e#�jT-�ڧab�����h�6l���]F5���mi�
E���z�݈WS�|���;I��u����ŧg�#��~O͒�=���W+K����zZ��������nf����{���;|Ȃ���5�~�u�Z�=�T�����t�q�h�9G"��\�r�4���a�f�5B�20��=?wZh�!j���Y����#A�d��+r:�������y
���!g�LS�8��0�Y��s��p2!�MB��y=,W�8?abZ�~]:�F����3���Nfo$�w�'f�������Y>Ade@{��'P]FD��sq�C�����U�i�p���3��bb��KWQ�6����1������Z���,6jPA���%^��=��gg;�z���P)N#c5B%$K����`V��^�aM	<�xL��0
�|N��,nY�3���5�!�r��i0�/RM"M氡��5?������W�5Z1����5�ԡ_��Mi��wJ:&�>C��:\ďN�����s�nE��y�=?ܨ.�!��N>���!��?��G�eҩA���|�������l�ZWS^�?���ly�©*��u�S�9V 0���npݐ���Ç�׫�����ୃ� yB���)���f���|g�O��S֐l�����/IcP�:�T�[.��)��ШO�'��:U�޶.z1�o��ï��@G���<~�-ws��V/O��/Q �B������A%֘����v�gYo���pĂt�X�=��t�F�A&�8ZFn;�Pp�O��Xʴu[��<�� @��P�У凾��"��嬯]ͽ9_���V��9����)e�D`"Y�T!�m��B�"���_#��C���w@�uP����Z��|X�PH�~P�c{��O2�7#��b7M��֭ru���� +�Ɋ�t�ҺZ�C���7�{�D��R��LO�o�2��2eły)(�y�M���P������LW��O��� ���\�F&_��U��zø$/@8�D�w�s+\�*�M��A2a��py,����A�ͭ�%�rJ=�xr�'�v��p�b%��@�d?n��H��{\�L%�j�˙�U�~Wq��r�ܸ ������Z�~�n8�7�W�ܡ`&�N\+��a��p�@�9 �Պjv�������de�>O?��\\�,�%xM�X�Z���q��W�oo�y�C<"@��d���F�"\���(��؄�U������7���.�y��2�M�1�_���Q���`8�@�
��t<c���:i�t��	M���?�*���?����l�<q���ׄl�! 	o�7��c�o3&9����[�B����hP�z�굓�j�h���$�%�6��=���R��c��kP��A���m[��F$��ߔX�ۉ�p�J�A�'�J�-I��f綺�:��cW��GN����	Є�74
7��#H��bF�39Ę�s�����uC��9jH��[G�p�ka?��pX�V}Ƒq�cw��sD�.�,]%�JbFj@��Ng"Y!��m�$�o���1��:�E��M�?��E�C�t|�t�+����xj�V��ū��&� �ZO�!�� ���7�` ���-n�����'�ߙG��O�_q�����6�s�Υ���������v�ǻU/����OPX���Z66��G+n�H#�s���Y-��s�g_���8Z�`Z��~��vkd,䔕E#������5��9^jP�k�)/g�<���T
�����'��OW����-7������?��3�a�����8^�Y,,,�3{.[L{"l'����qM�]��v�MK�|����K�����=���Rk6�ĨwI!�4����������Z7�t������BT�
gr7A;��8+�^ɓ +�Q��@.�	3��E�^..���W�����N.P)%��J��Cw�����7���� PQ����֕e�ߍ������̖�e�F�����/���T���~PQ=�茏���=8o�'h36Lz�B[G X�u'���P��c�Rw'�U������3�
���BaU"�k.ziiŏ�l�������끅9[;��IjZꔽ��\[׋vy�~x�L��@�ɨ�ja�fP����s��C� �v"��hbd8m�W�.���NP�N��R�*�Rccb�?�5[���-V�˿qyp��G�K�C�H�?����~,����N��#�2�	<�>���jl��Ikx0\�tC��j��赫x�8����O��sHGm���c��U%���#L��qķ�{���8Ku����|���ZU�.����%���{;Y/}�f2g�3��J����
	g��ߜ2�\�����1��r�E�Wj��e��jsҷ�UM�d�"�N�΃O)m!����1ޑB�3FC״@Bi����|j�7-�[��?�_�̇V��en2=�kr��"��`"��o����|~]�ןI����o�2	_8:3�盵Γ��Ha�Z$E�/fϷ�Vk�t��y���T��<|������TsE����"��������Ǵѕ�	H�w-�Mr��ڿ�~�l�Yx��><q�^f���2��B�w❉n*��Γ�d�v����C���U��t�7�k�n�H�GF�J�8�3_Cs��fT�=K[uQ[�֠i��͐=ߠ���0Rۤk��,TQ���G������S�nm���%��[0��+*��8t�J�-�s
YMg5d�۹��	������������m��N�Nh�� ����*��=OT�:�Y~�bE��Jt
hv�fy7�[{v��
%���N�G����ە�s�\W��n]��Z�z�*���o�p[hv��y�1�P,�+%/��-��m�o����v�)�lG�k�j��E'\,���C_|�$�Ți~�D�����9��c�5�ǽ��eR��E�de�iŃ ��n�嶍�SPQ�6�J�_�<��>p`������ڕb���jҟ�����fRRI˸����7�騢����C�42-��Y�]L�]6U�j�Di0&j;99e�Ań����-I=����'=q�����?��"Pad~�_�'8�6�^���V*��ΦO�Q%Y+D����<w�}$OW��|�kA��"�@�p�=A/��f�@�o���<�s7&�x'!�n\!� ����w����\'�/,{��/�]��۞��Z��]��f8�i�a�SF�2��0 �DtI�]a��|����:Xv��I�����7@�%���TaLÌ�FVK��tG��X�*�&�=�q�c�g��9�6�Lu��)��I573!���u=a5(��p��)2�G���J���ԃ�.+tsS����4��[�_tC��ڎ}�2��5/��u1ь4���7�4�aꯉMf��˨o�蹜���|�,-����ginI����l���XI�f�kIǓ�Ï뺴��1MN��:)�fE�_�\��/J3�Ծ$f% o�E��Q�q�ܜG����!�b�[έ�J���=�)-M!�)��&e���?�0ax�#�O0��ˎ�}�z���g,�ֽ� V�xWS�Y(�p:a������`/是:���(���I�g|Gofr�n�^�Q��v�fk\,N�G�3�W�;2R�X��\T�(r	�p��۝��-�J�j��M(�^?9-m�%{د+��窖Tuo�����9��G�~��*ce�풹@$)mB�r=e�ṵk�u�u���ik��ُQulm'�7^Kq���Pi��E�Z/�a�o�&ܦ��`YD�A[1��L��0h���m�s���Xg�U�U�:X�G퍓�c�����"��e��:��O�Eퟌ�l,�����a�����UN��{�>��N�Ғ�̚Y���(����$�{$�%WY�J���PJ����R/|��MB|�.v}7���ñ�b2��˲�v��	�?b�[�C���3_�h4��y�3��T}q׀'�he�B�nq�mJ�M�
��ĉ�4��Y��:���1g�y���t�������EM������-���uk�q�u�	�]�3����h(e�y������R��{�/���ڵs�m��O�����y�or-f�P8߈V��Oރuo4^@�ĳ��r,c/���K��"�t	���i]���;������'����3��W�Ӈ[aL��v�M���u��N~!�^\���_���6ۈ�Zx����2@�V�cg�}��bZQ��z&@�p>��_��B�|O�sH�R���l;���p���x.�[swM+L��p�Z~C׿�tL����o�E[��$�6-%�wNu�?�����~�j�����[�$4�&f0*�iI'/���f��x���XK�������Af�M^Z;~Gm���p��"�I$�JS�����gB��؃����fS:,,�?ւO��O��h�)}�C!3򥷏W0E�ep�H�Ԡv��
�Ȭ��D
��3��V�))��p̽�QS��,QL_�I;��f8`�%[­�J�E�K9&¥�8�Zo�h@�'''?U�`Zc����`��8I�h�zX�M�kw=��(�¾��NK�9�o2?==)��.��9� u#w�7�7�,[}�wo[f��2�7F�4�Or'I�4��L��M�첄l�N�/�����(
�먡9q�v^^þ�����s76|!B7�mB�P�<�`S���353�*.�:��E����K���	� ؔ�����tͼU�|�g����y�|"������S�wXi,�l�U�/�9��^�s�5�VRs�i��G�w�Ѫ,6�:/g�|/���IC�m����o�3�������O@-��%G��'�c;��ēW��[44��������$I���|
�d������^�P^��f[y��Y&Y3�.2��r>�!�
Ia��X��o����`$��,y7��@�\��oyY *�X�p�z_8&��I���TI�h�w��C^�ʌ�y}�A&���o�Gǈ��o�*��KKE�0U� ��=�����~���"og�qZf��<؏�{��5P���4�b3tB
����S����r9 ��Xn�쓑�C�֌�ե!��Gή��VFJ������9Y��6g�����U�/7H�X2!�I��e�Z>��3�;Or��&�i8�L�Yu9��|�� Q�Y!���g��@�D��}��;?�Ts��M��?
jf~a�싃����EQv{��eqGe2�I���gr��P+k�c�,��e��"�w�\.��p�ψ��0x��{�M� T�����=U?�M�E��h�}�&[)�D�5�k��]��^����t����J����ˮh��T�v�,��j�jU����[&ɣCdd�$w����"`AE���P>���z�S/w��^����h��X��5�)��TI�ϖ���g��G�4$��n�<NW�	7��j������>�9i�A��0��c���D����Q�XM�����jb���+i)��$U)oz�W�qG'߫�\V�`�C�ڽ�b�:(��S����}��_`n��n�}+�����/�A�Mg�vVq$�s�˪�JP�4 ��S�ۛs7ɳ�|��RM�N~\�l����kgO��ċ�#*<>}����(��~����!555a�b%��?Z�:���ǉ�swW��~���AMN������b���^iI�� ���]�y����O�gV׻���4��ͳ�u���u ��N�]Ś��a���������6O���Ff���jf%_S�m��gp��#:.�yq����1�sל~�$;E�����MW\�)n�4���@��瀆< ���/���!�ןx�K>J�mf'���&z�({Q�S3p%���nw!&�C�ڱ[�.=C]��
�'W�Md?�x�K^ڀ�0$ێ��=�w[����$����5��0,��k���_�3����rh�J�����M��n��cy���!��K��ƓYQ6sCM������o��.��BUH}X�l�ٴF+0��x(K`�7S#�� �â���c�Z�{8<�_K+Ƈ.�>QA�rXrÝ�o6&��?A��iܽd��0 ��W�Z��<��e([�}V�D���T��H�T�Rtn�캌s�?���,�2�Y�z������{���yh�o�M�)_�����my��<����{���W�lbj�]��%i���'9t����L�!�����AUmf{���{sP��j�_�sr��OE4�2�[�oc�6M|ť)₂�"欗M�.��=O���t!Q���	[}��G� ���/d��B"�;��=r���u\/?|��c���_Ƙ�¹u߁^RǗ͗�;"������&i�>G��gT������=���������\@b�K�?�?�ߒ�i=e���e�p[P�������{��gQ䨨��;�"�>�kR��_�fRQu��oGE>҃If��#�C�\��7=��z&"K>@'���<a���v�N�!ej��#���t��5�;Dҭ�N�����,�������c$2�X�($����  ��]���,��ɩ)�I�2�W��/�M���wn!���M����5�jyy�q�[,s��p2g"iTp#E���]�[}�%��T	l,D �M>²�Rq�(y�D�Gڮ-h7��e�z��G��Tܫ���g�mMrZ�~�:O��7�n�j%�L���Qԟ��Ti��R��~>v��X���L�,���W� R]��b�MIvr�涾���I9�ހa�Sn=Y�Rᇉ�+]�#�p�������m�("I�w����m�R_X�C��>�^[s*��B;����rʟj*r�����pS�mR�~v����O���	5f�����>����*���E���;�D�Œ"��t;u��c�ދ�oT
Wb�������+��䍚+0fe"�2�|ϊ��hV@�����aP^6"�|g=n�|��78��ۏ�ۦ��}�@֌��@4@Ig':R	6Z�ݩ��m+ف�{�"�-��0�"Ś�+�N�����-"G��m'"{]\w/`]����cy�7�����B�;�V��8��C���ͱ�Y�	L��EWgu�ݯ��Ԧ��DO����fϳaME����R� 2��}ϝ&�0��'�W�����¬i��S;���j����k��(�ݧVgncD��4<'�-���(_����*�\MBue�4��7���j�W�5|��F)�ԧՍ�lK��L���:��Kh�����6<bgVI;}%;�s햔T��l!���q���cU��X�^�.�XC"J�JL��F �ک�%g}?�vMML������5ۋXB�3M�*��#ղ-��T���t?ZC':}�����ڇ;��%z��4?g���gg�P�K�/�?�������J�ý�^�/��l5�[���&�r�]�%G�{�W��-�������� p��'nI$�A�Vw�΀��@qSL���T!=0N���ϕ�?u>�IgG�XFe���R� �L@E�L�+$��O*w��l�7)��C���֮�?v�Ϙ�N�=�JO>I�)��f2 �v��j��3�����DL�!�>n�&1�ïXZ��]z��kU�%;���l��}�t�yLdb�³S0~96b�4��Ԣr�bo���tu�A�JF���>A�%��|D`i��2�N7����G��Z��9��K�84%EoI^���Oן��M*�����-�=k�7V@��@/���m�lMt"�A��N+�#:��9ޅ��v�Z�eВݞ����䒞]gh���	�{����ϞL�x��/gU��L�o?_��aJR�Ta%N��2C()�h�H�h��YH���uM��)3��|��\dm���MC���c�V/�]m3J�\��H���A���G�~`��s��M�y�����iQ}��x�y.��OaIL'���_�{`L�c^�5\K�\E�~zbUK�J�o+->\4FUE:�'����/9�%њ�``P���"I~���@2�/{N�2x� gv���T� ����9�0��ߥ�Dj�
�VP����Z���ϛ�О;͟��\Vs��-�+H�|�2�1����� ��RXU�~�jg������|H_�k�<r�A�7�Q�'�i�g��}R��8���[#�]{w l�f<��T�~�>��W�=��4e�N�/mh�����V	؀�l��h6~�:���i��/�~L����U�P�2}����i:�!��3�cZ��2�G�5���0��$ٯ
a]��!ʭ"�,'C�񕃎-��ua0����H�/�=����Vb�{��d����b��fy	)�k��s4���?r�>hVj[2lv㙠`^�N�+&fl���4�a`���O�@�^�~.�M��9�	[��9�$]��(���j���1�8����wR�Aߚ�b�2=�m�_ ���_Z��?�lQ
E��,� $�G`�Z�Śx�un�	Q�:Febf�bf��	)��S��P5Ƹ*��m��)���_h��w� $�R>1����f����ⴤo����'�X]�$t�A���E`S�-� ��hl�,g��y<�Z�G,ݠB��?���R�.gM�QnR����$�D��e�����
b"_��?PK   ��W��Ƀk Jn /   images/8d0bbfdb-2662-4be1-b50d-e5d8de487479.png�w�&M�u۶m��m�vO۶m۶mLkڶ���q��w��9Oe�{#2*+�<./+�   +�CD��8  8��ڲn�3 :)�������4��K��� P��! � � ��� ��"���s� �� �
��/[����P �� �~�c��,  �������w �8#C࿳��+�T�?m��Bo��X�3@���p �F������'N�������4��������	�����V����Ǵ1q6 p���u�r�%����LOD�7��/���<����	���)����?�f�D����\��nnntn�tv�f􌜜��L�LL��N��N���8"&NF���v���\�y��������D&���d���H���������9[��/��<���[��W0.a;k;G%{#>6VVfV����S!o�nb�.bacb���>�����J�?7Uǿ��z/�!�����L�M��'�6p2�C�WB�I����?{;[[g'a;[S3G�����*�8�w��k>F�X����d0������w��/�_[�U����¥h�dg��K�������O�������.G#	[gG{�?�o���g�g��V�h���=b����b�ɗs��S��c���_�����>�.ￂ�)�������O��������>(��&>�(F)Q   	Aew�������c�])k�񩊪`4�P���*q�����u���m�Z�E�7R�����A]��_��R��o����� bڑݧp,Fw����������]_�vn�t�H�f#��yЙ�H��9��eq���M%�F�-��t� ��]9����?|s��z�M����B���0a-��Xʗk+��m��m0�Lܥ,2x˖��,����J��h����S�G�&{��d�ؚZ��S5�p��吀��`��F�@��s�*�Io�Ӗm�f�\6��4���T$��|�1N�u@�Li�����Z���/D{�Ĉk�uЦ�u��/B��.�M�R%ܖڕ��}��]��4�}�x3�3���>���U��tc�Ahc2zfbE�E�I�`��v$�D����3��x��p�C��K��0� ��o�6/�n�h8��S������Aj6��#��j���Wk�FG�H�h�y�����cHLd&�#Q��'���+D�ވ0�.;�I ������4G@����#��i�T�����S�y�-E�r�/���T4�tf��	��A��۠�@��S�Tӣ�U]Ƶ��h[������d&]�k�W�A2d�$P��� �1�k�U&��v�i�x� p�va�HD����=Ƀ�ֶ����	��y٫�����j&��O��.l�L֡Y��T寗�4w�a�röQ�v<!���_���˝�@sg���o�7S.����'BK�����qi��L���u��.�[Uvzrz���5n���jWl<bRϰ�
:�a� |�F۱s��y0�HjL�=��s&����˴6�����'7�W�Dw�(���5�$���JF;�c�"�ɏ�)B�,0U>v����o�vw|7[~m�~��*��#�ٝ��1��c�*�i"8��"��Yѿh�����V���s;��۞�SނMi�O�Ov���5y� ��* ^�?�����,�x�������GgN���c�:��Ԭ��F�fO��+�07�H/D�Y��S��ns��g)���~#� �q���>i饡�}E�������Z�����I<[��TS�� pĪ��~��PBh��}Y�-=��x:y_���a�8R���CU�oѠ�W3@:c�}��E�KG�7����|� �)��~�J\M��t���i��>8t���g��}a�N�y��P�ձUF� G��|e`�**�bV�~���
@����}��}�iԗ��s�WQ�MSb1������{�];gY�C^�H�t�(�~c�[����m�LJ��ۆ�J�`NE�΃��N�5Z/����3��8-Q���2;	gg���s�l����H������kxco�T���}��ҝL̊�d��ĵ�-k��D��W�<��E8�Lؐj�M2�w~U�ӆ�=Y���3v���|���CL`6�� ~�\�pE�$eݸcwL<s�m�3T�u�25����ZdX4Oq��嗭�O�w/feu@���1WQq	�lR�2�Sd�Z4�l�t�����E��+�;u '��3)j�D�uP'
���BЯZ|����G���o��uK��-�MY��+�vR�M�˫=��X��8�0b��u���4xkvX�z�Eo�m��S������A�|��0�&��P~wITk�`�s�7sV̉2�'���]��>:��V�1�4�W���**��� �-0S�z�E��4�¤�7[��O�iCU�A]ֳ�	����e�#.hL��i;����O��!7vX�՝���������mD���Q&&�K� hw�=t�*-_�}�	��r��6�2^#�y5��g�K�h�v�Ia�o��-��ߣ�Ts�J�Iu��?�{4zNU�hR��ʑ_q3}��>��CƖX����������Ƌ�T+0A�>���qXL�̟Τ��~<0�;�n�9q�Ó��9�"� �s�R�ۺ�%���v�q�5��Յ�A5��8��"��aMGBT T�Ӟ�5(�<6��)��T�5�15��9�l�����gՌ��Yr3o&�km9:�ʃ��}YI�𵫊Å�c�ۗo|�`���0[���X���&����Լt���y�&:�Z8��`�r��f2�y�J�x�A�E0[�6�#y7�ñ�L�l�m6�|N���ϸ�\��cE�E8`���l��{g��th�U�*@�g��Ue��gg�㋷��L�����́���-�dy8ˮ�믠C �1�oXd㑌���Rذ�� V �F$ �8�U�ڂ(�b�b����㿋��-�<��n����9��ہe�O��/k�6J�����bNA��Ԝ��-�?�;{~������6衪p�%/[�j����ɍ�S0<��M���up1ϧӛ�i�e���:�>�+�yc�(lJJ*QPu�N���f�:�9�����[�UES��)��aJsj<��s���VD5wge]�،�k��&9a˭��6�)��gv�r|Q��j��S7fۊN�j�@���t�8H�%���s�]�v{�wYқx�~萧~Y[ɢ-���:DM�OL7�<�'���
�	O��j���bj_�/y�2��}��%iV8.]�bK��
����q����慇:��=��O)U��!��3,��ˍmVB#j�p�.�;f�L
��}Wx�:'���1�7��\u�W"��[OS@E1�~�����:��(�l�pvwg��o<���}x9���,�8E�~l{�H��;TZt�=�#�[�Y0E�⩺����kH)���HP�G�6�fU�RRF��(�����_{E� ��w�ZU3Ap�Î}Ƈb��M-6)<u��}ɱ�-i�����T�j�4�M���T y���a��@��O[�oiOߟ:7���.�	`�t����]%��D�D�c@p����R���ļ�	��<9�V���*3�~��1�~I�x� ��E+:�f����������,7g���e GP&[acK��K6	�ԫ%�N��4` ѵ<cẕ��Z�J]�K9?�а�{;)DN��	�j������lJ��~C";7d�%�C�'�{�q�d"��D���S���( ~O蘏(�m1o
�����F��!d����Q�ľ��l���Ҧނ�q�Ul�����/��nȘI�ʠ��̿Ș��,���rk�鑌��SA��˰����rٰQ�Iڔq��jN�x��G�g�*~���H�K �����'�q
�ӫe	�x��ϭ�_"/��|�Y��V�x냵�m�%e��(z6Iȸb����{�we��e��)�v��)��=�w��k� *ᦨaC(�=�M�)*���"l����Պ*����<7�rs}杤�]�(�7�K�A�lSS�q�=���"��`�3���4@�0;e�
Ӆ"����/v�s#�$�5�����`p5s�5��Bxkʄ�C3T��b��}�`���,�y��>�(le-�2�4N�Y���0U�;ʓL�t�6��6�ŋ����Ŀht�����5�$`4 g�� ���OÏ���>��Q�I������u.�)���~x�w�O�.@��h|�`8�?�"jۜDH<A��.73����G	���1X�z s��=m;��y��Lu���U�.U1�B����njy��T2ӿ����������x��'���: �;e+l"�AII޴��ˊ^�SwiA�H�. ����ql�%��;�BtHL���`��T�0%�&t�,�t*"U�H�H���o������QX<�i!�ȴX���y@��o�͉�T�_��
=V|� �M{��$SLVg1�g����kwED������C�T��E{�fq��g��ݭWH�l&rG��)�{y��������a��4�8��x�jiV�̙t�)"e�� %ƣ[)X�8/CMu)�p��_��@��d��L��e"����E�%�����$�E��I-��\�^�d��m$�-��3�P�@A�{�C�J�E*I��آ��i�X4�oͻ��%�%7�7iL�saer� MKj����k��:�sHk_�L\���竵z�/����w��;��?h�vDB�7-�d�f�ʅ�)�;y��0_�a�Lm
�_ xY�xn����Y�]����;��b�v���H���?��U���g�&�e��[Y�YK���$ұq��>����v�)��o_X����J%6��ݣ`���)W�.�R�GjM7�J���qf���=�.8����hWC��c���qث���e��a��-���៱&�˙{ZK��;��X�ȯ�q�@���I^��r�>����%7Ho�▛R�������>��Q�?��9���_O�H�dmR��ᕱ�����X����8]�@�1�S�Ү����;�<�oᘼ��$���4��8��ɀ����4�v��LºH�ΐ��-�R��2T
��S��ɾL}�[2\ZW������ʋ�4���oq�ߒXI8h��I/+ko����I΢1#?Ygj'f�ˡt�E`�㾾WT�
6�(���;F��w�bm�$�׹n7��Z��u�w�Ecc#sΈ6��5 &W�E�&�i�/�;75�of"���#���&�s=�y����9(UO��Yk��C��Ь��� L�9:2�G$M��*tLsd�iiKl�/�An-hxd܏r %"ѼN�om%S	u+	7e�;#9�;�:���[��o�{�E�ew
�i,� ��W�(�3EE�2�VQ,y)My���0
8݉���u�?_�>��0������M�` �YI�BS�h�W�c����]�u�L)�ƕÎ�Z̷�_����6���BS��<���:t0$�x�U���Tb`y���g����`�l8M�բƸ�g�+�(�:?����RrD�M<\}���X�E��/��N�63��O{!a���ղ`\,��Utxc^ER�Ö	�;If��muurzwf×�)�K$H8Ŭn��,�Y�`����:N�*j��Ƙk�Q�h.D�sϫ�c-��w< �ή"���e�ܸu*L.��?F��J�����!.�}�<A�����.��ZL�;�W˰�c�g�<n��$�
��64��Ԣ���d`%�r��I��U@��Ǟ��W(���0�Z7"[�eи���d5]t�lh�䜅,x������	�{<�Q@|�p�P`�Z���[�~���J�M���`D}.��hT��n�F�T��.�8;o�6�5ܣ-�P*��~�g���	�����k?�3~Bܚ"���	��f��P������Q���D�ldmR�ZV�<O��e����.4:�����+ʻ!�uZ��;��]�:s�lJ��na��"]V�!�:���wCP��PZ���G_���:#�qi_>{	��H��Ů}E�y��~N(9U~պ�d�)^1]�'kH��4�͗������!��-Y�,'Gu�&��Fe�g9�T&Dn9,��hvy q�O@l?���C2ǔ�ﹴ��n�;JK��_�鎃���c3P �ԗ�j����9ðՋ"I����I֥-�`}�xYNs�J�S)����%�9�q�LHR�t���h��Ĵʽ��'�,��/���}��y�\��i��7#����-!,$Gq
��>��㎺E�0s�J����Z��#bT#YZ11*D�������g�y�rlfV�N��f.�V��5��w��IEZG�$�h�-�v�2�%��׎�fL�O�6�2��,��A2�Nt`�^&�����~&l��1�;N�"k"�-ZTb��<Z��kG��S�R/��f��5a�s+������IO	#�oLo�	�����ؽ����ƫ4�n���H�dBY���@�X �4_��*,z�SP��`y��z���t���<�J�\��TJ��U�7�k:���6/M��R=���w۠�Y��B	r8j1�_�D��:��u�%��nB�����i>���g�IP�r�F:#-*B�����4P@+��D\q���iж���oy�rEL�
��wc*y!���'������q�\eb�C0�+8C�=�|��p̵Vb$�!.���Pt�P�1,D'8<���3�h��?'���R%
w]Hز����)؟���.h���4êRPLzK-4�>��)|jD�"r��SY�iTS��P*�?��x���Y&��8I����	
�*B�\��3��q�]�!"��-͚�ڲiݳ!�6��f�>�s4���~_������F��-ܞ1�V�V��������u���p���)<�a^�?����<EB���&&���z8b~�G�j��W<A]|�}b;�1Ql�����9���e���6Z��!u�'Q$LOi�oELX>�9�&F�Llr��11���d��I`�L���C��.5F,U@���ѳ>I'f�&|�����
L��t�J���ّ�L���|�<OpE D�Q����Ǜ:�p���A��,�(�C��L��ل�4�|� /��9]ҭ#�+Q��Gm�U@�s��O�+zB!���
�0��j��x>�XĜ��J�Пy�=�ΙU�W�;�LM����<��R�f�����x f ۈf&q�,��O����/�<����-�bb�����/�Z߃[��VXq+,��4�i��c�[Jl����}d=4��^���y�"w��T:�ǽ�׏B���Lf���uP�S_��%B(�8 )I �+Ǚ��!�u����ʹ���o_�s���.�4�(���J�4�������a���F�V��&
�\H���:�q{uD�
�pE��٘�ʳ�&_q˷�z���qH�Ys�/ ��O���2�ˑs�uY�"Pp&p������1qwzp�b{EX��?���Pqq�r�R���V �J=�S~+��3�i0$���VXv]��~A�)���^�s�_���q�i:����߸�Swe������D*ao1~�]��K����<��!�'�e��
XT3`�aNx�B������.VzC�Ԩ*�p�KC�߬A�]d�Gt6���[�d�3�eC�`쭌uz� ׃���`��aG,�K'���>V��!7��B���3�t�}�2Я@R�n͉I�6��g_��W{S�9��v
��8�F��k��XG���< ��h�	 ��"�s���pK�����o|��>~(�;Y~%�Mŀp��R�=i��HcazNP�bI`4H����	���	�)w�|���q[�]��d���p:a�q�؏i��\��X��:����{/�`݆��h� /�b@��4��:�\Y�����{��q�>�\`O��r�XE�R-6�i�yJ��^��0��l�ߺʽ��t��e��P��c�E�4̽�TD�Ad���g��p*���}@�v寋��!wiG�2%u)�*�4�>�v��b�J䣐�T6�!	���@��d��*,��j�9�o�M "`�T�n�v 6^y�K���h,�v�,�.���J��?a�[��װ��gix����[��h�.kb�O<|̐��n�9.u�kG�9&o�ށ����g�*��>{f�'<̈́)��*M��q#LG�#��H͡��|W��5^�>1����| ���- ���_m"�r�����.�W���SKm�����?��O}S��v5,}H�wP�~Ύ��ix �<u|$�7�͈g��n�:_�N�BH�F%���iU�n<X�C7R�������g"990b6�.bYy+��o�H+hi��|�`Ȩ���Z�q.�~y�` �?�~~7Gб|zg�݌?B���n��x���[AT9��a��S�����rK��W��ww��T�6�[�Pqϓu⾵͑��ƿ4��2�+	�^�SI�.�o<H��2���@��p��	@��(�������l������tt�jxц�Z���Y�`�C�6Y�V����(͖�B�x�M�:��������c.Z/|C����D��I#ȯ��9�u����y�l3��/#/�ꆛ �QLh�r�i��ϲ���)E��B-F;2��^T	5�;��n�|�bˉ�	�uYk����X_�����0;�$�?��T�#�7��vfvR�NeӼ�����R����Z���D����g"�4𵟑{g�u9�ZŅ��76$������}dV$z�@>�U���:'��S�l@�Q)��3y�"�c��v�q?9����B��՞�D���LӈAǯe�S�z2�s*ޥ%Es���x���G'<&��+`A]��$��K�26c�j���p��$e���8�2��+������)@/~:f��9?�f�,0��A,��}<�LA��W����ζ�'7t?����Zq�^>�5n˽ ;/�C҆_���(�V2�9
鬲�wO�I���cy*S��G�:#�Q9~ ������<�f#M������T�=B8�,�/���Hz	�0���O�M�x�w�ܲ�3�u0N{Ӈb��+���
no�P��(��m�`��C���,��x�����mq+�/�/��',��noZ&�M�d�2�]4�7p�w�ib����b�A�꙰FR����P�ę�x�tcO�#s��ʳ��=�N�j����r�;�egSb����+�C��lp2��}���‧6��C����4N6�Hb��'3z�E}�(S�Yv6ԩ,�,���q�?}U/_�y4����2枥}���zH��ʏw�$�(��ݘ��Hh�G��{u�eQ|s�#gd�)����L�nP��4.A\A���pF��_�Oى���
��W"x~�ۅvASiQ#��uIc��>���������'En��F�;���rL�% �L�$�ukK��۟�c'ûSnp�h����{kg2[qU��_2j���-��-�D��2��a�n�2O��ї:XG�C��a�����?�~����"�.�k�!�"ֵ\[�݃�	s>w��2L��j��n��فy8����K�KZ%y��i�^H@��d=FUfIc1,]�M��$�d~Ձ7)4�� �I�6�Mc�Ҫ&@�E>�=����"i{^p�b������]_����U�I>�)���/z<��e �s��f�r&�V��l}�����C	�l��U�%;G�䤏��$Z,�k�fݶ�R�S��\!`^LH�z�B�n���b�8@:oF��!�,I�5� �xi��9�P��.h,e��
&�������\Yh�E/���`�A�K�q�*���*�qRO�o�5��V��2#�$�C�\�b�J��q!� �2ن��I�°�%��vܰP�7�nd��/��S�3+�b�5:��)n��k�,u���V��[����}���|��ɟ��v�r*,_4<T����� V !����G�?�%����7�j&�����=�'�<�\P�@/��aUg4�P!r-�Ɍ�+'��/��k��'Q��{�Rל�OL�iHȔ���Q5�B���-�R���7�����-㶉bհ���7�ɬj�a��P�R�(��Z�`�n��_�������i@	U_�$Գ���p~�O���AANh�e,�[X�g�yp�����p������H��%G+�h-ݸ��k	�hސR��/:B�`�9�\����Ć
�A�����E"�S1I�M�~h�g�H@�q>gd2��xǇ���	�4�LJ(=��7�&�}4�5⅂�^�$w	���k5�]k+�K�fh/�;/�ѵ�I7��Uӯ��z����g�<�{3�m�DƏ����0��9'g�.���t��`�HΤ1��S 2Y<��c�9b0�)�C�������k�Fa�O�_b�VM�f�P�2cҤ_Mt#Br��ڸt�),u�DC!��&櫥�,&Ώ,�ʕ����0�n� h����zQ:l #��ά�38 a@p)��`1�S��+������3G^8%H�� �� b̎��[�e"�\�)T^�dâQǣ�n���3�lR+�M��޻n}@ �Iy�"���P�l�Ǡ/����<�&AXF)nyV��@�}�1s��nŃc��V�aj��-�b�s�|�@�Aӈ�E��P�0K艸���S0��
jX���˸�}�d�<�C~�Ș:��tɋ�0�.��c�F#2�ڎ�,����,���	�E�v\ƨS��(#�:#�!\J��
8~���[6��:�8ɘ��?O�M|�E�^����Qou&3{��Qߡ�ώ�@�5#Ic>f�T��1nv��m]Edq]X�؃c�:�Zkw��ѓkg���}�u�~�a\�ab�KB:�(:��=�j����l���;2���7��r��e��5������R����$��.��T$������*j��������{��8����?7��W[}�aۓ��
�8(z[�A�D�����^:bf0�y��)�;�+1΢�O�S��s����Pw$~Sʕ��N}�\�]�@�vZO�!��V��ɤV\����1ŵ��B:��Nڨ�җV�~��>�Uh�M�+=�����+��U��q.��JBQ� �g�ϺEX�ˆI�&�U�*�0b�r鰏q��)?2��Y%̗\�TIG���y���^�y�� -0�P��3\��Q9K-��WC5]S��+�0���z�!z�xli�V�4�.�6�������T�ڏ�S�FmP�
� /�$���a��L�}|<+Q��<,a�K�ݥr)dE!6&błYCM�WX��;d�C��MOMՀ�2QR�ܲ_\�[��c�d& ��O��GJ>UO�����P�>gA�X�_��3HV��菓��*��>�4&��$�ߏ^&�\_jiFe�M[H��ss���"z�3���R�+����6�������`�@X�P_Om/9��@* �	:"���@�aՀ��YC�P�=�,�Mj;�&$��b?�cFr�L�ۈ�ڝ��K1�P(��vN���9�M�C���5Gw�O����%Y7]��GA�~��;+��K�;��s�SH�hėZ6�t��iS��0�e�eS��o�_�ʻ����E*$Q�O���)�H n�!������D<����E���<Gk��=�τi�c���M$ޖw]�co�B���!Q��م�����Oϟ
�pLĕL<�iD&G�����qq�7���76w���P�)Fe�t�I�0T�� -����H�O������}��ZP��ה�%���'���=x�W����k�.�e��#-(܌4I�������	�.Y8�
��<-4������B#��.)�4��t���Z�V�S���kr
%�h�6Z�)�~�qc8�"S8�~�;h�4�d�>������
$r`8�~	.b�P~�ӯ׸]&hA2��%A�Yˇ��U�a=���49IT��;4�3�{��EK9�_�zc��a��{'�X6ԁ��5���*�ߑdXN�X�ש�������L��A��Q�j�P�8�R�0R:���%?E�d�k!�
B��
���}�D���ZP�07#�+�u2�Iu�g\5y�e�'�y��qn1&7�A8P�7�x7���� ���&ز�d��nR͊#*]i����B� �.J~\����R7�bNTd�rL��A�j��"��\�Z<d� ��\�ua��3叚�x�@e ��΁�Ĕ� �͚B�@+'e�y��=+`q'�����{�~�p�7⧇8��F�(#���j0|_q����P��\�wɆbQLx�Vf�i9|C���Q����3���p���`f\bs�R�L���+)Ґ!�&�e����	�@5�Ұ9Y��fa�	�P����
��
�tUx!:K@�K)��$G�S��&����O"��G������@p1U��X�4�9*���W��YRf��%H0e^���2'g�P��A���@���@���2*E�t+�ְ��g��Z,T��h>)�N�I��v����
�H>��;B��mG��:�s��n���l6S9��.�$��!��=�-��𽽛�(�("H��H���|����xѾo>��%"�.#a�UĿ>�'�Xe�\T@�ve������&��8������j��D`|)���dF���D����,-aRٟ��=RQ�c�:*��ߎyL����U��XW��8��Q(���z�lRK)�����w�� �K6,�Y3V�U�:|��(>|%���G�T?{��0�pGuo/l0�<l��Oc�*/�yp�rnؙbǼ]!�ɠ"�Ŋ�912'�$
�E���.ҟ�_�^��yhXL�߯�ɗ���z�\u�<�86�n.?}��BeH@-#,�5�Z���)�{6��-��A��\���%����W��(h9�A��LGuбy/�3C�0w����8��V��|�^]R�l)�Gi9o�M`hR���}}�4ځ�)�fũd/�l��H~��d��F�W�:�� ����H� L����<e�i���ݣ�'�GK�����Z�2���w�A�j���H�kS��p;G��V�ePk�&��:6��Kh��$�`+�	�4C~oė�uJEvYL::�52 ���S4�R�hܩU�cY��ꏘ�u))�G��u��*V%��x�z�Z2�1q�z�(�k���Y-�:K�1�~�u�e�����_�?LeJ���]���(����@|Q��Y5sZ�C��3�Eo#�/BG��B��9�tN�2�`6���XFB))�@_".��Es�Ē��e�803Ǝ6��[��W����Q��)N�s�oS%� 2R񖠌D �],�v�H0Y���@2n��1�:�J��E��6�ׇ��^`��7��>F�6��&��hx��Ql� �9��}A;V� m��Z��P�e��D�G,�-��Q;�tn&Ez�ґ$��'�!�>^|���P����ٞ�Mgކ�j䝊��9k�Ƞ�T��(G���1�r��n�-l��IC�h������~BI�VYJ�[�C��pcd��_[-803#�^w���h��4����?�0�g�Q�Βu��U���u�es�%<m	i>x���D�Y"]��mO�����l|[G(�%���� �6��h(���X�6�&	��ج<	��&hu=���0�m�W�T�Ӊ���[��&.��a(䂨X����Wr� w"`'�Ga닒�Sl�g�64�i�O������H檚*��8v�V����r^@a;��J�
 ��0<�@[|�¶�`,US<�Zi�#�3LK�O- �k�j�y�r���X��\������w�Ŷ8\����І�A��G95�W,s�������7�J�5l��\5�����U "����(����[v��	�Q'\�8�L�vwV~��,ش)0�.a�z����8�[B�ʖ�ޥ�qc���)�bx�w��1mT�,�WG�\��Ύ�!�i8�~��#��aG�1!P)�}�Ul�\���r�G��2�y��KdjP`��e�3bI�IB�0`��7FhW���%S���$��wFWx�������U��l�����	��<$�eF�Ȕ��-aIY�%ֽnԞƖ��sD��@&��������lC�cY�U������)ELuE��D�4��A � -���ag0��BJT��F�3x0�ts' ����9O��Юp>BG��e4�+�/��@�����	˟���i	�n����4���Iz��ܼb��Z@e�n@j_>�� ���%=���5~dI��$FP����D� ��U,��:Q���y�(�R-Z��^B���b��Hcn�	����,<v�UX+�K�J`C���Ә����2����i�9l�yP�]5S�[9@4��ma����(�	0���|�V��1EW��\�;?U�Aa�"�_�Ed#�f
�Z�M��W��N#��)^w\��?t��^�8�"���f�+�r���Cś7��ʑ�ƻ�+O��4��$D䭔Uk,=Z�sd!X�"^�wEۛu��t<>����t(� �T�r�:j��C�t���Qg�n�0Rv��e�|qQ47U���`�yB��C`xE.-&�B$��,��|�\F09Xd�ir�.�J �|ޢ��>S[Z��"9L�WF������VR`ݮ�ͺ"�`�Y�{��V+�Ϲk�Q0�
���2r���/x��-L�Q�z@LJ��G_�CT�*�Z�� �oQ�z��{v�����dF�iM�EW3�{U.�WE`ƣ�<��X���O���>!UHZH���yB����_,V%P+R#��f�^�o�_�_z�ω���UiA�[e��/��`�����^�����!���S���֒�)���c��Ȣ���26v��U��>���3���O{��UJ�hVm ��4@e��+Q���GBӓ~�z5�M=.>�U*��΃��0<�WItfk�J�������9�sw���?��4R��Eƹ"�8��"T%%;��W��XG��O�2�s�������yt���~��v��uk�}�78[��Ѩ�W�f2odغ������5FSI�*=`�
*���ȳ{��K�fͥ�ʺ�7�����z�q�X��赆L�G��Ç	W1l-f�Ʉ���=Q�:7�Ѳ&_H�2�ڳ=e
��/SJVL��'�Xp�w�NNl"2����p���I�K�n�"�	�p��ۃ��Yڼ�C;�Y���70�hp�ғ���$�{^*md��t��LY���P�6`����D#�0�ȑ<ks[-t�5���|^-�i[�4�?���A�r��4{��`�y��ۢ��xb�)>>1����"��zN �tø�8��s������>���$�J(�1u�^ꉟZ����Ox�p/LL���C����;z�@��6�+h���0=ZF�>�+1X�&��H%$~�A�R1�w`�h�0+���a(C��G:�<��C�q��a��r:��FZ���q�SȺ��c��Q�i����1���uZ����S�4|p�����C���5��i$yfķW�{=
j����JJ3�2i���ȕk6�{ZF�eR�_�J�xC��F>tM��BR��r�!RZ�q"HBaZ,]l	�br�)X!$�FaպHW����n���7�wfmoM�}��%_w��cQ����,�*��I�ip�Q#�0�A�����We��/�b�p��=䯃���f�F#-AW6и8�x!�xW��ո���4���,FT����H���+G&L-�QF� .j-:�2Î����Ϝ��"��s�%[ۊ�������,�:�A/{�m�Ü�0�ۛ3]>o���:�7
�6xq�2%6*����rn�-�>Y�{9?�RV�u�.����>o�:#�����y�}��dV�tx�;��z�쾹����:_�z�y���P��Φ=�?�`����ҴDG#x�b:��[�͢�����fേR������]�ظ5(��ݬǔ��"�5�K"����Ld��v�{�v/�&
��h�M_F�e!�l&��B�Z"�j>'�����%�����}�#xэB�ze���K�<
��#���f�ܿ�J�)$A�av��9O�a	Gx"0�%F��D���m�ޕ�[��9��θVF�ݔS{�T.W��n�l����������w��ԫ��1�7����lE�II��R�cJ�YᴂUg�����u�_����s��8�6����F��>�:��:%B��lB�~�mm3�	��X��4j�͜�@2�%��i/]��RE\k@ C��9��2}�aU�5�v����uJ;�(��1����!@޿!Q�4b�� c�˦p)�[��&>�3 �����@����5�=@Kd�s�\��]��K�q ��Y���֫)s�K�2�
Ŧ0VZ^f3Q�<L!�#���&brBшBR��c����c�~1��dD\�,�P�N��P����24���^Q���@nƮ�`�#�d����'��e��I��l�2q��!�Ԩ�3� ��&s��bN�ۮ�̦�G�ẜl�t*�WLv+^"p�1:E߁��0����?�s9�H)��݀�.9ݺ�@��i��Ԣ�aH�'�P�0�  ���@S]�4�l�"5d7:K��g�����.R���2����� �=��I�S�`�1����KM V-��p%F���B�&�8{z)0.�x�:-�_��ƈ���
��r�9O�Ap���Ƨ���,gY�q@�S��/b�3KI�l����,3�.��u@^��iO(3�PR�dd!"d-Tz��3aU�܁l-LJ�=�W��i��ΘM.�  @ IDAT�	eH��m��fR<���(�:vL%��������&M"��=�[�0�5� ��9���j!�U����J�Y��+"�D�i~��Ur�G9!%I����ܚTDь"��A&l1��U>�@�z��U���XT}�*V$���[zL���]�c@��cC�R�K�r�ƫ��4=e�Ë)mNj�!t�T�$b ���(�@�u����\���+j�1G�����7��Ѹ��!��]df�$k5~�m���(<4}m��k�����[:�x��S�V9%<�I�&VВOy���B��`�(�j�@4.Ԭ���#T����1����J3Ù��Ɍ�u�h�Mԅ{�A�@<$P��=j����E+Q��EoL����6Lņၐ�;������܂�a��ɍ��K�����v����g��r�HU��@4uM��r�R1�r�!vC�T�]�~�D8C ����W"DR<A6rr���z�R�tޢ"<�����ek���-�yW�=�z��(����3�Qx��A�%h�A��ݬ #�>HIߑO���җe���T4:V]�"�|v����ά�R�O�����j�gC��R[m�*!t�Y��M�Ӛ? ,��2Ϋ9�N�a �U�f`�t�R�j����|�oJ�#�n��L��/f�i��w��*��ʮǥfQ�f~��&3�$e��ōZ�ka��n��4�dfj�J��)x"�+�F~�/�FӖVJM�>Q��dCݫ�<ZEҥT�p�@�P��լ�*e�_g��p\H����*9��#O0ʃd���O�+E*�r�_��X�OƆ�f{e�PT�B*i/��OpPEJV(��&m}��(U��4�AA1�V�����.0�R3��v�"��� �L��`+V����#f�M�Qj���)��bd�~���z8}�I����m¡CB����x�����g�e�����_ݙ&�4hv�e6��4���+�Kd���3 (pUD猢&	��yr�G�A@f�q�b����l��N/t}��C���ʰ�p��CY4n� M����҉4)8�������(}=	 2���q�
�<>�Э�`���Ue3��=�+H�w�� �@i��2�В3Lػ�ޗ�X8�4p�2�@sp�LQ(���!9�-�qA�R�h��m/��$5�"�)�'����C��jZj��z��,-�XH���;������L	S�;�����Eϒ�^�&�ȟJ�@Ϫ%�
��ؤ8���n����]�f�,"^��J�VX=��U�>T�J�)t��m!a�����Y�vT�B���8r��=Q@������0O��9�.�Ç�l��R��TB �c�&��\%Q� q4���W!(�/���3��
�٢��yf�)3 ;���	�8o
�$��d���4+VR��a���U�Vk����tb���ı�\ys\T�\-'�G��.%�LRS,ϴ�a1`�*FJ��Z���o0� <xd���GE� �y!�55 Y���C�ҨP�jM�l'������gsL,Q"b.�L,��	[?�27Fnt̪���mɓ��n��1�8���i�*	5ߏ��}��dC,5��#<���+�[�`�*��*Ma#Q��оEB˄!�v�F��G�����3���'I��� ���UH���x�����_����.&��@���|ụBH+�Ok��3��dgԽS���,j������@9!�C~uMt*��YD�, �yӋ��\((EE"j����pf&\Ql 2zhu��\��Z�:'XWd��M����k^"b sMfP@�*-��Siq���,�p[�O
�ӫpl���R�AåN�,�b��u&�j�a{U я��l���F�R��j��'�%@�h���I�PN�\����-��.#�1�w�[��>��A���T0uB��A�Q��B-��O�Y�$��N�i��u.E#%�;(@��H��t&W�iVt�<^d<�C�t�����o
5��8�W�if�ꔌ���V����*�;)��D�@�e�\���)�\��
t?hJ�(�a��"�ͽ��i��N���v&�q�/�\~ ϻ��r�Q=� �M���5��N�����~[!��%^�a�܎ݫ�]��Ya��9<�#S������Gz��`�L�	�LA�j�{��=�i���ɨ�Z�J$W���t'�(E�~�3�X������i� 7��<�&��
����{�<Y�^�@A����7��r`��|{���̔�<ɛ&y�3��$����'�-g�ٶ]�m�����}FȞ��c��H��o�1O{p}��8y�N&�A�
o9Gd�f�B�ث�� 2]����gH��1U�����H$*�p�� (U?ƾ�!$\o�{�J#�B��9 �@��H�IKE8�Q~9ȡA ��/��f<����웨��o�L9Z�| ����6�a�!V��*�P�����\u���eX����I��P���,o�'RP�� ��x���W����٨��7��d��D�Ҵ�"�眓S�d�����/Tg�/�f��g�����VQ@�iqY)�Hn(c#�0g�W���q�-M��u���PP�g ��#$�f|�m"��V3�&�m	|i�|E^��1���O����C��Ox�0D8�Nj�1��W&�p�\k��Y QCl=�-�����HIx���;49�~���G�=y�e�a�G�A��żA����e�ݵh?)N�tD:5���m�B�0��8����sY��!���7_�
�&���b�W��ntXy���n��1h�ԎQJ:��e�9$B��G�{ХӔ
bۍ�̴������h%[�^4"�ͥr����:΅����j�zqs�r����&�v�ctj��P���0a���? �#�3��X+�"�b�ɵ�
��cն���D'y �߯x|_�?�!����~��_��ן��_��_����w���ڏc(+K(ND��V�9�[����CzHH���N���ֺb�1:���a�ش����~3�K�,o���x�L��C=_|��W�߾X�ܞ�s<��?x7�xw��J&�Ծi��,�v��qU7�Ÿ1��y��Թ����7���b0x����1[#�w��jO�T������7t�` �;�7+�y]�������m3��b1�600��-V /�Mx'�fr���ۏ=�\ �Gˮ�"�*`tj��X���HA�09�RH�M�w��������뗯(�?����_����o~�/����}�b��l�3���1o���Z�F�Fe�a*ft�mn:�z�D�b��"��"���A5k'����t��������^��n���XF�v�Ӿ��Y,�(��)CB9o��l1��z�m8�/f�ռ?�.���7����m��j�QL�(y�����Y+č^�Jt�|ouV��m�r��l�s����:[&:����1�fh�����g�J��\���\-�R�T= �q���\��I'
���m*&?�����_�����~�����JN]���DԨ�������(_����� s͊ｲ�j�\���x7�ŋ��Z�헃���js�K�H�}��ro�i���ƺ�#'Q����y��v��o�����d2���$G�գ�`��jAW7��M�b�6Μ�A�K�-���M�Zh&�b����>���w*P��c1yI��Ƭ,��I�ȹF?�#�0���ͤrfZ��N<}Q��gѴ��e��,���}���W�/���O?]��Β�+e��.�k���れ.��)�X�_ac���f���ӆ�������R`��`���
u�K�\B��i��o,Z^�g!qX���g?�����z8��o_�z�o�c5��gӳ�Z�tFw�fƯ(w:ώG�i�Q��׻!��'@��+��zT�����c��zn#C�ySq�Q3�Qq4���
�h~���(Z���յo���=�o?y}/ͮ�[��Y_~��W�^����GA�h���1!0��H��ѩ$��L�j�p��r
^���o�����1����r���Q���vK�v���!��PV,�u���T�]������g�٢��łN���C�Mo��*��u�V��\[�f�z0�q�����F�j��pu1��G��#�Tz�1`�%G�T�u�k�.:Q�
�׫��Q�Gۻ�*!_.�
�
Mi!�E�0Id���ޑy|�a�����0�]l���y]&M�xa�t��o��M� JK�=�R�'!$G��Y�M�Wk�ǍXW�x����q�
/�k�L��%4��K`���o����p>��Do:���%��>�{��wu��;��� ��^i<�qO���C�,?�"���@����죆�*V�r�+[`
��*@FQ�L�8K"�ڃ��b���]3�Q�w���h�|x�S�x�����@5Ѣy0�ͻ�$��UQ��O��������AFŬ�z�D5�m�������j����lm��Q�]r�2u�v�BT��N����u��o`'_s���k&*��8[�! g�^-w�+*�7��`R<N�s	~��'���yJ��{���SEu��+�Ǥ�}�arV:G�,F&�n�� ��*R%t|P��i�H������y�Ĵ�-�6��GgO0�֬����<�w}�n��qdT�m��
���5�]�Y+B��0�J�	=���XMڡ���O-�H�:/��V��i��9:;�]>�/��ٹ�	� $�֫m1�!�җ6��UF��0J<lY�.y�� )�2�:��0�_���x>��H��M=�O�B�J�-�f%&��㢜#�Z�)�\2#5�lt�&�����X��kI���w��a���u@z���I)��R�p�Zs$xб恨(��O�]t$h���}�i��9�JV�n�N��y����U�U�\�	D�4h橴NǱ�(0&8����l���n=���ө��N�矠�zNc�h�z����ٛ���rp��v�[ķ�%������1�����$|C[Vg����`-�����L��]�g��DCͭ�T��5@*X�@j0.&~裘���.�>�S3~��/��/�Gdj���f��F}:܅'��k�u2���~KU;���g�}��w�iUV���T�8M��B�S	�n��v_���X�*O��>��ԉU����ϭǥ�DN����TU39��d��͛��3���ء'
� K������*�ΐ�d2ը��#`� c�!���bS����)�e=،��]��p�rM9/��'�d�,G�,�������9���F5X�v������+�)�k�p�K�3�W^R��a�E�7t�ScB!��?e�p��S�ȏ�~y�������_����p\]��{z?X
�2
�P�W��ǿ������i��o(͛�����[�We^�g���@�`��s�Z�;�9���)�AF֬%kN�Pe\��Jl�7A	��P_�V7g�S��h9�e������g��6��e����d�z��2��ۖϞ<���y���3�X��3�w�������o!5?Y�|M#��P"ʬ9�!u8,g)Xs���Z�C߻@{F�"	��^����k*x>[>y���'�2P-G���,Y��H8|F��r4����֋��vvy���W/n�u����]�j�ܳ�)b��M�Y��̳��$����2}_����T8F e�_jI�M�Uq�I2	%ξ�*�""*�s_/�p�5>;���z?����cl&�s/�UU���wg����1OA�nv�5˫�,g���?L���a����\���$�&��� ���z�LI�E���1�x-*�AK�"-�?�LqR�裏��[��Ʌ?��w��WW�)����;.�8~��G��������+�i֜�%c�,�d!/:8����w'������J���o2���@��ӛ0�R!�� c2CQ�Pp�ycVM�&2��*:�,�Sv�Ў_Oow�s>����B�&�cN�*8+����^dd;G2F�����¯fJ�lD��i��y��m�SꇞP-�R���7L˨�i �<�XӢ�%� �t�Jȶ�h����w�����W_}���t�\�ub*�����]�᪌dA!/`ξ1L��^�F52���ٛ�gO?���Q�h�a�T;����/(j�����ڂ.��e�\����yek�l��|̆tƹ#��@v��(�OB3���-��,�
�KEXrS�j����55��T�N��E�:@BX�O/[&�'\���kb::uE/:��3Ɏ	-�6�3��n� %g?�336�$\[�Q���A�
6�d��B`��<x-�{�}|�q0�)?���޲�������N�U���Ti�B�MB�,�?����xrqs5�3B�������v!q��r�����a�4`�k���#bF󇸼�1uƭi�\,�K-ޙ��Å�S7*��	i����Y3,m�r���n��/�����r��`8z�a��B����v�xUr�6��A�Ho^��{1�Ю���t^�}8���j����Q�� c���{G:/�G�H�Y�H��|���˿\,��^���okg *�$�x=D�P��VT}����v��t=������� ��{}�L����НT��g���"�#	�OO�$����Yj�`ͷ#b��R��8_�
�� �"`���fW!��b�f�����������)rc?�x2�ѧ�~�������E/��7�]|��%/̧| �7��h>�}���b���c�?����x�:����zģU���5lߕ�?mG�s�Q�h�bnXqBk#���h]c�s����[rg��iE0�-}{ TiT�]�56�l8���_�I���pzu�ւ��'D4b(Z"����bžE�ի0���'�0�i�`q\9�C�����d،�L�;a�8C�!tN�l����t������)��T��;�iWHB���%1Z�F/�Y��k�����v0�����^q��7?��ǃs������˿�}���8��ɨz�x�oV�:Ⱦ#����ľ Z��`��0�W�
=tn�L�5K��K�0բ>�4��Pސ�I.Ԑ��hN*�M&K3nT~b�mm�ٛ�.��~u1:sqUY�ι
���^D	�?�-W)!L����˗gZ�s"��+6 &�b�.kX3{L���&#J���S58��'���@�����T�;�=�#~d|\�������~�u$z`�)m�}�6��dEM"H
�XL���1�~���L�,��W[m�� ���j"�U� ��9[T�g��cv'c�2��c~̡o���|~�U��bԍ�=D���h0
��:�0ĉX��ďl>pk��lf>�5��~ղfщ�U�㗉Ix�ظ�"9Pu��-�, �l�B  F�(��|�ᕧ{Q
�����+,2���,�����#@1�K5 �%9�����4
A��==6G) sڙ(x�:
9����c:�K��eƍF��KjC̢<�	�Ț^A�yٹJ�Z�D5��~��%7���g��N�*@Bl*g���m�����8�R�ԏ�~�q~���V,h�K�0����!|*Y)�6�c�Ѝ�bB�d����f�s�Ы5��- 8:om+���`��t��i hO�N2���MCG� 8�!��b���_id߈N|ih��O��&�A�r�Zo�!�=�"��qAF�Y��a��P`62P54In�uT��@ FR6��;���8B]��rѣ�!� *�9�~�+�`Ν�7�x�u��פ*,/)�C<���[+M���,`OuC4�<&��	��G�Z����rN<;_�:`�ƒ?��s�zmy�ɀR02�����h*�XB����>��\R��]���	�L��M3 �R���Ӛ��	�t�0SB�a����uAlOM� k��5w���C�{�yw�%5''l���d����0m"�b��P�5�,�Q�U-�}���b(n�tNvk��*���8����nzkM�����+o��BV��� �s��eo�tmQ��Ͼ6q�����M�:��Ctt:|��r���7/���A�0��d~�
C6{4�d�O���	X��8F���;����|-�Ć9ŏ��&X�6�1iQR3�������	H]8`����v�f�����/�o7�>c������AB�
hv5׽;���ܸb Cެ����_!i�=$C�ʎ`#�G�����.��_��;���@ֆ��/��:!�{s���~�T#V����nX٥� Sw���-�Q%�{�!�Au��x]q�.n��zW.��Ag�W��rw�WQ ���QazGИ��4T�ž��	W�=XpR_#�b嵸��R�O���6c>`�d<�C�H#s� �p���͛9�Y�*�7�uG���SVL�J�2~�#�n�D\�H������;�}_ךu��!#�3��f�&*�����,�E�=wlD���EQV��|��ף>������П�-���*w���:Z��Q�7�S|�*d�^�E-�8,V�	��l��ͮ� �úx��/��d9�Y3-w���U��-�^Y[0�2$hT�0�
1���R 2;�z��PL}�N�����	�6��lX�����;2���N�ɬ�7�qx;��?��z�3�9ɇ������c��G�<&���%c$C_�_��W��lt�$bEG�t�����U30d�B��`����{�jSLjDј��/8���!-��*�!�+W��Gϟ�|��0��|�h�f�O]�d�E]��dʃ? �͂�u7��P��E���|8z3|����M�
+mD7-'�Y���n�=>(�ͱvɯPz��k�̚1#c�v�}Ɔ�,f�XM'+��V��JB�h�M&2B��U.T-/��t���G��/���_��^�]�}sɊ���E:1�6���b��w�t��7�X��Q<J%�n.Jn�Q������Y���l��b0BQ`�\W�OzSN����˨h�d@��(0A�A���B�Ԫ�_���S�>-~2Ҽ�o����O�(�>�0����7��3����)�N5�����V�H�*!�t3���9o�m6|y�&t�׵iw�c7�+ˌ�b��_}��_��7��Y���9���)"��7[I{�u���KK�K�ހ�*(�A�⺲�[潴G���++�!��Ζ.2s����ِ��尙?+6�_�_ߎ?���з��ycK	>s�t�R���X��,���ޟn�ݛ�t�ڊo	��]�X����o�Ͼd�����)J�15A�h�&��y�A�JHT9�+�4��K���Ps6$ab2I��k�������ӧ&1R�=EôF��SP�����l���]Q��!��Շ���Yxm���V��o�a���q���s��%�'��p�a�PǄ�hb&"�#�UI��@�Sp�%�:Ts��/�	��ɀk-?Q�-�f<lΛy�zy�-��ޜ)i��<�G�?"��[nF��n1^��i7���U���,n��|Wgت��Ӵ�B�n�H��4��ړ�e
�2�'�LH*ؚ���_�eh|Rƶ+T���RJ(�:��2pB&��e�	� {V�ua�_-��$���#�`^��3*�F��x��1���U��	/���N�"�� Ӗu�&d����S^=4>���
��Q�p��^��E>9^6�I4��j�~����G�Y�w��B���y��r�@5��7���n��Yjf�2tWTQ�F���sr�J�G����t�[<�@�e�Fg[m����r��([{����ՊWj.u�����0�i�I�=� O1I�߬�t-W���>(��۸U��9j�T�Q+���W�A!�1��Q�K�|�7��N��������:u������.�H(�<�6b���}? �kJ�"�J�lTn}�`ӛ�{����5��g��ٖ�y1�v�Т5}B۫�[*��9Ӌ\�gK"���AU������k�0�@߉OB¡l�-�j�C��Dc	��3�=�j�:^�p�A��8pk�7 �L��Ql����*8�z��})V�c����TB�@_������{�=�鈞��+0%Qv�A�ۭ|�����c�8��l<V�m�x�5�ڵig�&�"���? ;������/Y֦&��VWKV���܂�����jc
G&�U�:�N-�˃4M�Q��É Ea��?
��ĩ�����[�	�G8� �0C��G�ם].�9?ԢMu��!1�c�թ���	4E[�!2v㤾ɧ���2���0*�5�H�YW؟�Y=%�V��r���Dn�襰�9�9V�a_��vUo�7kFWC^����p��qM
�����#���pLO��I�E�i�Uo6�ގ��XnXQ���bǬ)U�Q6��r_=�"�3S{����v����Ƃ�E�&ՉS��]�=� �F�Ț9T�H�U�a}9V�� �}��G2a=����'
%r6�O��an�4> ���g�#�/2���-N�Ⱥ�1���V
9Ӥ�������i�[��Up`��ɠ8������f2���V�A��ď�d�Θ���T *����7���;^�D��ť�
:S�K�\������ %`�`�aj9��	*���pf ���@��8�r<��IԽ�<�����#����焃o�@�LO�1"��*��|���1���ZP�!
�O�m"8x�?�NK�!M�j��x��3�W��XY�
g֪"�8�=��(L�5� +��'��K��Y�0:�9�3�ғ��k7����C2ˣ�bL��K���V�S6��`��o���?��fs��a0��m��YF�p<1�5�N�͢�Ex6;�"`���k(�w��Lp��q�ˬ%zL%l�x�"�X]V�2���'ܙ~"�d��D�q �y(G�A3�Av�!�ب��\���=;?g ��w�}��G��wyy�L2���&F1D�ь�FnV����/�,kv�z��|�����M����dB�4��0��&�ge�>+�?�޳I�$[�K�3K4�h��sG�ݹ��K#͖�����\Ҍ�/ܫ�6{g{zD�t���J�)"��{<"*KBU5z���._?������YvXv��2�*�]H�*��� �*�[��3Ք��a�}��i�tL^8��x����>�}TT5�.Φ���,\Q��aQcJS�1-��LX��^@�Ҋ��_���;0q&�ł�&# tP�~�D����9�7H� �QW�(�"Bb�ý,f�����od�Eh���2�& Yj$lý���m(]��N�Ra=۬��I�4���-�<���Y"CC��d�~3�Ũa¬��)�!��r)��{e�$�ǽB8ΰ<)�Y8	\��XG�F�ՒD4y�.B�Q,r������{��2a �C�i�)�)�P�bd��0�c�+�y�b"����f�+k긙)�C��M�%�t��R�Hh`�'�J��2�-^��b�(��&|)��P�S<ܯr�=�j}��d���/x��TS�ʥ����z�xQ��@G�R9_��wЮ���?� �)t�bȏ˼�R��b`�1\�|b����$X��+�y%�+K�v+_*������hW\������pZ��E���ع|8�3x��#+(�E��z�bV����@&JM.�������af�����`M�&�(��ԝq�!�o !��V%�U��IŮ����$ֻ�V%�E�ÏH�A�	Ґ�Q�K1W�+�\)�sk�.�A�/y�>r����}.���eE�I�}ˈ�ee� ?/�����bL8�o�b��in=���lB����|�����r\����'O�^��#8#޼y�T�<���K;sͯ#����V}�6��IP��Y�G1��(ל�\P�TŝC8G�Qq~�1�KK����xJr 2&=��G�F0h�RS)���
�of��pA�@Y�S���8F1м��#~�q���QF7�x*�������h&
~!8JbA:	�TBXc`~�0������û����Qn6��0�5��hپ��5k�~�30��7�9�x����*T���s����nk��}뽷9��)�bM��w������!��Tf�ٺp�����t5��רk��8��49,�_��0<�c���'�2��U2v����;��P� �P��z�2M%2��ք���;�Q���-�KY�^Kb��Q���$�����A�O�p��Nv�����=�ϕ�"x�-G�M�C˘��F�N�<}��߅����X�kk+��j�}��vWV��ɀt�5�Z��p͋�� ���u,8`:�V+�ݽn�����:�^��fu	'�֯
�ޯqͫέn!~���%.e�p�\Ǝ]թ��9�5y����f�-����a�zn�a߇�Zm���Ũ�B���f��2�'��q����Y`ⅢRYNQ��;qƤ�`"9w'�)T��!��18�������8���zp��ёK>=0ji�V��F<%݀���0�Lw�=���)K�Q� �1'ƿ���҅��F�݁�u;{(En޸�������J�7������?����Z]]aY/T�g;���Րy�l�7¼w#��=�-Q���<�3�<����5��ű'�����h{|��WF�!��5��؟�?�H	�̘��$D���9���Y��������=M$r�*�H�~2e�d�&�πB�����|�8�-?�ɏ�S^:XW\.����z�f�es�D'!��-��rh	C���������y0��#�,K��R��|��ѣ�_ކ��|�ֵk7���ڭvk��9Ǝ��p�����(����g�%S�t�������A8a�:�=WV�x��bR���D���pf�.Ģ�U�r�l�.�8����9�(+��Y���� z�=1k�=�Ti�44b?�&�h/���X�}0��*�ǡ!S3�G���2ė�''��|���y��e���O�"<Jʁ�#����%�ihi����kB\#�/qA#/Q�dWY�1�&�D�(ص�m`�ȡ\('�ͤ�S�;����_�q��/߻{瓏���]Y]��/~��q����v��z����_�܍����6�;����G�Z^Z�m���W��u�V��C����{�����,���ɣV��'c�ln��w��
x�����%b�0Jd�SE	�aG���PC����>�2�Ķ��F]�8�s/T�QR�x�.i�����:c���������nĭ�*-��G�kPX�-���L���3Kj��:=�եH�&�4�/�K]-tw�u�씒�HB�!p|���\/bX������D��Y���8�����ʕk�W�7���V���c9�ғ'Oww�?��G�4��<PU.T���۷���k^�e$6���F�r���?�iss]S)�X�7�$N�C&jɟ�eVO��3�RG*��N�ָB�����dG;�;	�-֟F���R�?(����PŹ*���r#�h#u�`�喃�)"P,zʍ��i7��W4P2�b( $�H�n+Ǉ� fCHQ�	K�ռj	�K����(��z�Ǻ��̑��~c��rC�|��!�
��ĲQ�����9й~�*�[[������j�!���/���kׯ�:���^����t��o���Gz�e!�����*���E��BA%����t����Y�s���M�0*#� �cjR=ҁ@qi`*�eŗBܖ���cV+�P���~��B��������-P��	��$'P�1��JƤ4��վ�75���I[*��P;�920���K(K�Z�X^ZZ���E~P�1+�����B�ϔ�hT��9��� MG'e�����kW1F�yÓ��{�Ŧ�I��v�	Ѕ�
��&��%�D,'+���sw<��d.�.��9�"D�w��=��u
T � DB5o4c)�k݌���U��V;�<)�s�����	X��
2�Q�t��%���x,����)�pīyvf�e�ϔ8� �\K Q�|�L�t��WWV�� 2Ɨ�b6Z�Js6�e�WwH`!ԭxk��ںy�-2�����z��.��Ֆ+�A����ݻwa�K���y=�:?͊2��X�ݷ
	����e�?,��l�E�@�0(z�1�f��6��U�<���̘���^�����I�Є�h��\�l>�ڏ�0�H FKiX�u���V^VBfZ�����EDl��
�����-&��"8K�GY�h�P}�r�Z.]�tz��Θ>*�9��݁t�Ke� �L�|K�0ZYY����Q���Wk5$I ıZ�S𺱹�lj�����0��B8{��j���9�˿V�E����8#�6I�HevӸ��nT��"����S����rx;��*���-���},��`ڝ̿��æ�&ô9:���%2���+:���}�%h�B��Ϭ�J�ń`������y���A�V
�i�_��Sc�j�a��kj�P�\�p����'�~���F�	D{�4���˗�2�����f�P`�� b�^�p��G˫��9Ȟ�
�R�k6�0��D��Y���s� �Q�� ���_�ŷN�K<�bb�A���h���U���;]�)P�i^vd}�>���;����f���=x��'��L���la�h�RM�J��x`��R{��N�MG�s���V^vM�b&u}c�Kn\������	|��n`X���eY^��p8*ײ�V��J����sl,�6�!�ۺf�����j�b�� ���z���k׮�T�p�f�	�쥊d�$G΍��.ȹ��a�9L�_����@#����ؾ���W�\���8r��CwF(�@�l�j��/�����]��p̓8'�,���\e36&�0�H�M��\�%������rX �����f{��������M;�7;}��]ޥ2�VYf��4/	�	VUQ,�y��$�,si�i�-v�1��Z�ճ�_�u�������Z!�����r6]Jϊ3�7�cvh��+,<q=�F'�m2O߰"XRQ�;��*�"=r%�ն<���<�nT@�袰���z�-�099t��� �rz�`����?�9p<���[NΑ��`����b�/|.�]T�F��x�B4�����at�1D)eW��h��ԟ�;�t��w<��ޣ�a�Y��7���k�JRز��ʗY�j!kc'�3Ht�-I�2����?M��T�/���/��������s�څ���ܰ7XCW���Ҭ�o�A�*L̝Zs�. ��Y���`m�����/���N�d�o�q�v�{T��" 0�+6 ��Қ�L��ߺ�Py���?�����m���Y�8�j���<�&'W��1�)ƙ�%�:�@�T�����ی�d���sgA���ǭ�R��3������k���^z������)�"��0H�y�B̓)@`�E�+�C�]�x�=2s��ػ"�f=��v<91��}��2J�z�k~�\�S�Pּ
x�L��z�igo�����Xdg�O2So	<a ��j�`��V`2��Z ��0$�K��̌G�8�����v⸛�3���3�`Wu��L��֮���o��Cf؃�����y����]k6��k��_8c=1\H<ύ`�lE�^K����8DQ}��|�D��8h�3 @�sF-�x���D�~输�Y�M�(Q ,�{P����XW���\y8Ɍ�^������~�x�';�v�XZ�2���G�vC��l"�-Ӓ@�;�HL<fAEa�FS�xht4f;  _e���<sD��	Teo�a��a����!�LF����ӭͥ߾ru�v���f}	�0��˞>T�c����]�ft\��n��<�&ciL�Po(_ ������d�]M�D�F�jU���f�a��[�?�{�m�w��i3�Y����������ʗء�8���1<B��ݟ�����ݠ�%�Dt��y�IS�������� [���b4�n���Kf�S�jl��ݾ�^����Z������h��GAG�)���y��+��ḯ�)�5��Փ��T<��Xs��� �?�>����?��;j���Ti�d҆U�W`�� ��=qCN��� D�G�&M����w5^�Θw!mt��+�Yvt�X��i  @ IDAT�]��Ű����J�\��$���֚��f��Z������n��^��zQ��cZQ%
:����F�bqF�������3�븊��I���6�qΣK�}��vw�O���� ����5'�G+���P�06Ly��~����Z��������aPY�{� _��Qp���d�ꋸ0�Q�d���Wt"k<���XA��x`3�Q5U�X��Kb�"�H�C㏪�f���c�[?]���0�h���������˫��w�4]�s�Ҥd�}�w�(��?��_���GwFggC��eIx�?\x2�����5�l�u���P��U��DIDKh
�MP8�4���S�=?3),�����o�����˽�R�Xf=L��	 
��%�#B��d��K�p�!!��ֱ�] ���dneA\Q�L�	�������E�������K��2��eۨ����e����Nj&1|�3������?�M�޾��5��o���L�_�������R�4`F�-�"�`Ӑ�%��ā����F���Jhɜj~�/����":'�pB�ݥ[÷�(9?�%ѝ~"��~�˘�A��N�ֲ4-KMҼ�PI�R)��#����n�����y���`']fʃLn�Ύ�h !�x+y����$g�`�dc0�p�%tÃA]�#5�ߺ�ʊA�C�:�f��8��$t�f4�5<�)�"�nʁ	&r�Ƴ -`JK�t�w���$��~���|(�NL>cq(B�u����vf'����@���-�w�%#��-����l1�=�($�Z�RN��r|�G,p��|��;[�����}��l>������4_�6�%���.��u.9F��Q�!8;~0ØF����Dw\��!���Q �����/�N'��JERr�!gE����Q��\sS[��o��jM(��ad;~�/����h����f�T�4'�N�<V��i�d��B��y2�xJM�T5���x�n��A��Q�Ɍ	_�A�Z\]k��Ͽ}�_>���v�I{�����!��R�&ѐ�-d�6�9(��4��j��4��F�"R���A ��X7��q��"X�G1�D�4U�)B�0�n�Ѳ�ʷ@H��sL-�D��}	�1W���_
:[ww��Χ���7?y�Bu%Sd�2ϳ��!��fl��JB5d��:�@A�������\�g2��8�.ΕH��Q����K�C���ȉ)���$<�2�^�E���xЙN��|��mo��׏>��ν��k�����_���X��>��������!��9���ɩ�9Ag�X���B�R��Y^�.ɜ��Ԗ<�d�L)(T��f��A�w��H�͌��B0�5�!Z�0�����	jJ�!̥SO�ݺWg�u����퇻��7?��'�V'�ɴ��(i�k��q9�3Ve��)ˬ��g�Ho�ɘH��$�F!i/}�?z��|u(��l@v(�3�t�I�Taj��J�l�Y���ýO�~����C�L�gI;�-�B�4�t�k����k⼴����C䘦��q3+3�٘��r/��,#� |$�A�hG������1�V��1[�A%dS��@2%�Q9;Ul�SI�dI�]`�q�0󪕕;�g�;��\}4���<���a����k�4"S�w�����d�Ϩ0�Y��4K����p��w��<��i�Rc���1e(M��F3��ɝ0ԋf��
�.�A�P�@f@��|�
}�Ӈ.MY;&8���, x��]�A�`�%�(�E��Ω��T&�ɉ-Ce��NuR�n;�	��l�	�m9ôf��+����o�z�j6����w��Y<�b%�b5!}I#E$XT���qt�{	*�����n�����~�>a�{��j�������������o�>J�4^�
��RǴ������ٳ���#���,�f���B�IdL8+	hZ,ZD{b���<���{���9�]r��%:$&J<@M��"{�|t�z6H�=6���*�:<�h�
�YR�3U(3���%e�.*�]}�����ߙ�}����8I�$�)�c���a�6r�!\'o4<d� �):D�M�/�a�EH@Ms�r�?���$ �3�^jG�%-��6\��a��#����4�n���gJ�ڽ�{������z����]�'36)�Z 2��?�G��y�g=$��3�R}�g��l��E���`e��"[$+^����m� �d��u�Z?�1��Zn���R�ZLX5��h%6�P�Z��%4� qE/S���Ϊ�|�; o�z��n�\oT+��0������Rh�+���@ˌ^�X�˦�9|UN�*�'��~~c����:�#���UVB�1�=3H��$s��b躐U����,L��X/�_x>��/mup����7�'9�R�S.�1k(b'��������n�8ʰU4lH�` �(���� 1dzy&5�w17�F�jw�:�2 ý���	R����i����z��Β�P u�J!��36���f'a��b 7�S�?�Λ��C�б�W��}ӵ�W�F�Ɛ64���B��!�䉉-�B3͂l���>��q�P���{sc�����r��*�n�T7���ța�@e���7	2W^;I�*����c?�`����w�����|�UX�1�3�$����7Q�Z����Y���h*1����S�t0��S�Ǫu�3S7���-=�9Q�A�,�t�L�0>̰�&F�!{L�!���`�Qe>��*��2�V�;�| ġ� Cdu��/ϧ�^��Yr%�c��h�0ԏ��H�i�|V�066�zw��=�>��A�\Y_��\j��Y���ތ�	:߯������A��G���SIvn��7i ���g��ro��ow�i��kW�^-���ߊ_@��fl�'s8QB���.�ifg����(��{�b�=��F欀��4,��=t�6���
ᴸ�-�l����5���w�ZX*{�^PJ�a���ʹ�ߍF�.WV.
ӄ�R�m9��ao؂��Zc�N�G�s��(�QQDLO���v-],7*��#�ӻ�֗s�Q����.�z�2X0�O�X�¹�"�y(�J͵ܑ��d��YB�( �C�k�C=I��C�;��@��Cb�>I��7���� d��f���n������ �@��*�dG�e�\�����B�~�YЬ��\�U+m�����|<��IN��|)��'�i�I���O�m�[ݞW_a�+��vw��7.������dg9.S@�K)���,`�y����L���/�z�������O<�2k6��a2n�ƞ�5j/�ra��-�����Bz\J���;�PVԴ�X�z��e2��0�:��hS�6�`8���u�\�X�+ ��̣�O~���{AvT���U���� �D�(�3�$����V�6I�s����������^\�Z7��Y^{���4�ƣFƤ�\�����<lN�����vz$�%���N!7}ks��_���F���#
�Tvt��n��7�hf*5R��)=l�,�I��dP�:�!�ȅ��>%	2̂��kT�{��y=wyٻT[J�Y�t�/��
�����ޡ��3J�Hk?�a����S-���UK_=�����]�^��S~�r*���<7��1���I�{�	���^�� �����f��FjZ//����\�'a�1 �0x���j>����>�*�������!����K��Zj��bI��5�uĪ�(�F�\:5`�Iu�_wg���N�kщ�� -r �+�Zd@�(@�5B��K�y��w)n�\��_}s�2[����G�HcFH$ �s���_���&�$M���9�LB�bRԁh����K62���^��۷?{������u�J�� � d���B�i�,~X5��s?��Բ ���O��i�НɎ�E��2��;U�����,�j+�u/�~�g�K!�}�U����J��Z��w
W�8��ڊ�
(��I[:�?�\���>.�H��I�^Vf�����"�P����/��,����&.��G�f*�v�����<�r���U<�"������%V�r������3={uJ�@
aDтb+����w�ů�k�P=��CCC	Ui��&R&"T�g�����G����|�����^�U7=*����kc��!�X�|V-�W ���hBm<I���=��%�@�?�o7;�_X�\�~���q��bZ�8�5$M�΁���0�VM]�\fr��8��w]i��5ܨ� ��U��3{�>~/�p4%%��>̎��4�:�f}�Rmi)u�+w�n͘�`�:�#f��N����#����s�͔�De42A��t&�Ѭ�Z���(�������f&�I��]��\+�%�Y�EwY&.%4��A�Ys�B==n����ϣ@�N�E�rp~A��~I���jzB����,�������� [��k�|YJK<�L��b{	h��1	a Jq¸�ȹ�!%R;ў��h�i��K����P:h�����1�ӈ�!j�

 ����h�4��"�S Ų���5��5a�B��B��cy:�API�A�-۴7�|���K���"i��o~���N��3+���v/UH�k�����kq[s���s'�I�(�"�\���|A���sϩ�$WKP+̸ ��(2��y���o�u|�|�����~hB�Ԓ��D�P�~6T�R�,��#V\�J���[;#f�1+�1���y3�E�U:������۞�Ы��vX̢� �\��k��C¹�;*1׎��<��b�����w�0H��`�Q��z,��g�a,�M~��-��2[��������4����:	a$�_�s�ǋENuK�%RB}1���`o|��� �f���W�yeG�Ao���4&�0S��P ^Ԃv�C�:�"�{x!���l0sS�;�Q|��"1Cg�"N�h@�w#y^BQ/�DiO�����g��E�`�����"�H0S�������z����_z�<*'�ǻ�ol�pV��q� ��x^(?���e���d��ٱ��p?	$���2��~����qg"��0�j�R��l}z��X�XM��]l<�i�y����H`�~�H����zr�Q�<�t��^_v�Z+@{�K0=���*W|%����W*d6W��j���K�A�M�`�qp����b��d���.�T,��O��+4�272�Ij2
���xoCM#`�8�=�#��7�~(��8[g+���ޣ��&Y��u��I"31j��ً�iR"�G\��h�/��߿�א�1(�P��|Y��N��>���a�9�hz�؄�Წ�Q�|�W��.�8�TN���0��~C��jn0�|�#�+@F�
�� J��r.�q+��+(��)�U�RŉC�PN k����PA�����#��"�/�N["��(�k9z�x��?#'&�#Vp�)/=�|q�Q��2Y�(�Jqwrv��	�=	god� L;�Yyˇ�<�O�~���n{Vn�]��;~�SPC����0	���0C��`�ŦI4"C�! va�^�����F4 o"I�9��Mˑ��xW�x
Ȓ��M/իHV���=.�'��F�)��ᣟ��bѧ�0�����(P�	����"�<|��>�M���4���y��Du�耾�����(G�{3Y9�0�3Z��p�x�熩��V;�N���d��ȱ��2#x%$�L[����f������W���������kEe`^�K�fb9&���'$�t8�DY�R��,5c.�R2S �!A'+ y�Cwwf��dl��V��Z�B�E��43]�t(�6�[f7ơ�����D�� WČ�M�љ��7�w�rkČz:���r��	�{(�WYBE
�N�ȡ�.�ˉ�?��X�f�=�'d_�߾}7HW���2�Q�¾Xz(;4�=̹`��Ŏ@��虣:���`�8F?�+��4���M�+<z�ci�?���7F�w�� ݇�u���':�PN�A�Y3��� ��y`�#�~����`#S^@ݲ�<�k7֮��x���t�e�9Y�"sX����l+���TQ�Ug3v�-�S(M�=A�bF�L��u��՝0��o<��҆�Wt/A�����\x����a�)m���������.��97�8��˗��q���H�I{E�h�a�+��wIA�i5Gl��Q0佂YR�T@Md��P �-����錱0D�� ��=ߵ{.lH{JYP�<���աL������,<�ɀnAyC����1�#$=K���%ÏFĂ�#U��ۺ�#�I�8�:��'$6�Nf��d3˷������;�w6��ta<�Cz�o����E+�y,���.�{s��+Ř<](�tz��<��,E!���`�,��PJi��U ~�>�0q�p絟8+?W(�l7'�V��l:��lf����^/��z�R��"jN�Gg
yA�<@�kП0k~�K�2�ʐx��k:�]�-�U �&8@��!��N��\1��ϒ�i�s��$�1�������>t����hRl,#u,�f��:�~lQ�X���=����~�B�Q����;���3WG�Ъ_�S�R�4'��������~�Ɉ�p��g
��7�D���r���1�_� ds���y%x��3��1h�-�!O ��>¢����c��"���f�Kjb��9u�c�� �ꁪp
<�@�$F����0�W�J�{$��#w���+��Z�hIx��o[����0S���/�?��.ե�}��	d���HAN����g_5cC���n���s�/�vL�h��*`J?��4;O�;���TR�����&�z�!�6���ŵ�,{.C�z]��IIm&�J�� ��1<�H�C܅��_~�4O�v�����J�҉I�b�\�R��JD�k����-�A��'����l>,Vv��G�.�"Co0���8�E���Z��w����g�%�_d/����Lpf�#��p��G��Q��D-g=\5�*HQ2�UM���ɏ����f~�F�2n�s��9��;����z�"~Y?4��uyG��)	a$&�J����"BdD�ۇ"ѣ8���iҖ�l`��#��\@���,�����!��SP���fۣ��fw��rJuL���c�X^�H�O��̓;%��<"����R�?�W0�r�>��N�GE�I��.%�I������n����� i/Y[�CU�r0򷙆a>��AW����ť�)�HI���<��e��%?�����m1,T,}B��-���:D����P����҅C��7�L (CN@�a\[�}�B&������V�����.�	�P7�o�_ꡢ�I�/B�����;�D܉�F��\A��e���I������~�B��c8��k�@y`L�k� _�A�h��2��I��+�p��C��R���`<��!�s�
J亷�"��m�o+w�����L���s�[#e̓ (��E��$I���`y��E����e��3��Q8�JP1���C�����O[&44�I�A*��9��eL+{�Y�R�=Տ��?�<��!
1���K���N)-���2z:�½�N���sC�NZ�f��Yu>Р�����cN�u��g]i�g5��|y��6�C�t(!�R��W��~����Xт�3�>C���`N�8�',���7�XQ�����2��?iUʵ�`�4��h�5�P9ό���ܢ�Mz�kL�j��>[�i=�|�9���BVw5[Z]�o
��I�p��^�)��;��0�� �+�<���Xw���:�"\Ψk>��`�2g�M��b�ڌYQ45,0%�{�Z��l�c�U����K8�
Ust��$�v)$�2L��xm��Ћ�E��hϕ�Q	ʺ����V��@%r(�ˉ�]��P]J��#���!(\�\��5��"��WdJ(�A�]�D�"p�%���������ZY�����V�Ʀ+)����n��l��,�<��	I:��W.O?���?t`L��:*b�Q�1YS&m5_�{�D�h�2vP쪭�e
�>V��(�t��*����|V�
aVQm��.��F�'�����0xʧ�ms�k��(Q%���3�^����J`W���U�`2�d-���h���� F�D&�eX�`�ƽK9�͂��Qa�Z��8��*
�je��:����e�ƛ��Mp���U<,��j
O���aY�!�T܋�������ݐb�NI;x�bh��Q�C4��,��l5�}��������H��:.΃)�|���ɯ�IR��v�O��0V
��8f�i�E����@��Y(8�Y�S�\���l��:����?�1�M*z(JQd�~"-�R)e[R�Gc�� �(1,P��&��s�h',��)6���PrX��"��XB� h0Gʔ������]��y'I�����l�1f�P2�&K�m�A�SSY(HR�8�D\�o��_*��o�+唗��Q����%�4M�m�A�#�T��(Qu�:�4C��ʺ&*��RI>џ�^�R�'M�Sh	�C�1Z��L4���9�!�ɷ����?�3��	[������/��6[�|a��4,P,�6g$��x蓵]kjL�dp(Y�X&{  �C�1�u��h9gl��卌sB�I0�W��2���1��t�"LS�:�Pu���$dKFN���K��������IU�-rg�#m0��Y��&����b[���`��w��t��4��$$�Xg�6��+	��
aqD4�-{Z{8��lM ��|D����x�yG�W��L�B����
�-)�śc�!�mi�
h��:}�.a�6ʚb��\�}E�\�e�;֣c0�.�\i�}}l*��)�YO ���9E�g��u�D��'I��~T/U����>��ݽ�/��} %Q=��X⩂�R��I Շ�I�����Mi����B�ov�#p�L+%�-qgG��!1iV1�b(e��Q���<�:�;�j��$��M8����ᘭ���)����G-�8���UW;���:��ͱ�
��^ik{w�E�w|Xx��O�y�1�;9w'�:�<��s.a�c��&0�E�~|�����C�M4Z(��͌�8���!���P2��z%z�3�.�_Q���GQH!����ȟa�!�6�$mGr�7	�?rt�. =ċ�vz��tV/�C,�4��[S�FY����X��ҁmc�*l��G�o��7�r	���I���3�'��H��"PsMHa�Ɉi*K�	�k��#���?���:��c?;�!��c��2t�'�t�J���T3��w�B�I�7�
(�<�Bn��+�m4#ɨ�9���Hqh�� %��0&��a+k*%�����H�C:�����j0B8�m�����+*f$�q��}�qL�Z �+��b�F�4j�FGÂfz����ZD�c)�C�����&���_��Ra�i` \D���
�b�~�p�o�=5��M��ڊi2AX%�
i1�Ô,d))�*��ܤf�[H:pda&e�d�ǲA_�̈I���ȡd�T�FTn�u�'���5��'}�ǃ��W_�&D�r"��Gc�J89}�&�����$Et+�q�XN�6�Aa��0�sI�@O|�x���wܩ��cC��`���v-������WH�&axUI���[�"�L�0����޲w�'��K��s�Z(M��"���1N\�k�Ea\�]�\<WbL���׺����&���謆��y���
��jH���=��K,/��6x�^�ʫ~FWAH����� q(�����H�Q��|>��)-ݝ�F���M�h�bT���sc�,����h�%޴�b<aU�$�R5V����W؉�^������%&��#uo8�V|T� qz��Q[`�D��Q%7����ȕdDO5]��"vj��?�Q&ES����0��l�>	Ԕ%~l�($kٱ�F��D�W4̎�MX|b7^��^>Z<wq�V�/��$�q���|�8\ŹԮ�a2I��uiZ£�s��P���J���" c�(.�'by�!ڋؠZ�6����al��D������I,�,�_؎% AoBg�%�%ɧj�{S9tR�d4&�,!���M�P�t:˘��ӐP��YZw�(5��ٞO�h!�M�)��'Rb5�	�~���)cl��)!�p���}�����nRi�'��PzD��ģ��P�y��m��6*��`(4qa��������l�d)2#� aE�A.��>�ZP��CH�\. T�;�Ɍ���q���5�.��b0Omo�2 d(ad���=,���9��Phr�ʧgVY��)="�cz�k�9`q�\t<W�ς��oÝ�e��g��� �!�N�<͔�'���~�G����~�;���.�ߎ��n�8W��c��?�3�WzG�'j����QC;��|/��(]���o9��u��V>�C�����Y�AdS�0�#�E�?@A|�5�-��u4E`���(U;�@��?'�MRp'iuN���e�Vs�0>f�J}Z����<6}:��G�;����;�(b�,U"?x�]V��A=R�Nʳn-rE�:8�"[.�	j��8D@�yMVe��ޠ�j0/$q[�W��D �\+�j���2ģ���%�˰/~A��Ώ9�il0�ex-��ː�����x��1�[�ˋ�^��q��d�v8��Y)�6����ؕ�cn�z+)rrr��/ﱱ��ɀ�s���idkAX��U�ӰHm������7Yzd�x��\�h�Y2�����J�&)9J�e\j%`K���/�B��.`D��Ϝ={a,���+��Y����Dv�������A�4��8��N�6ˑS�NŅ� F9X�"i@_��`���?�rE��(��2v�2R�G;^�yf�!gd��u���q 8OP����RL*�f�qtj���8���\�C�	AF���L��L0�4*ZD	ñ�(=�.��.�i��V�R�{�����c��h|�fX� D������5�X3�j��,��I@a��y�''"i��(�=Ƥit[~k(��(�N�@������pՕ��h*�;�wo�X��זPbd��J��v���\�9X9]m�S(=�)���b�{	����'��\C�l(+��K��hɇ��wQX~�da��P0��lgIQ(*[�%�[�3���#6�Xj00����w�iR��/-U��` 	�(	6�"$����N�<�H�;ZƢÉ�.����*9�ä"��dM]�uA�Ľ~屵
Cl�X	������'b��;�iZ����ϾV�	�r8W���c+��a�7<�i��x����9�:e�h�s���kJK����@�yX��O�%U�Z-�;���4�vƻu�0��;�!!�@�J���v :�֤�l'ˌ��NT?����M����|)�D�R�tfIo�d���i霔�+�?�dhZ���R���Q�T+�Q0����-sQi5�G͢��N
(�^�}�5Ja�wf�lp)��P:�O�O��)u�Dw%��y���7QA�a� ��A�	��:)��`4�a�(@� �d]_	ɪ���^PS)��&�1� >Q���q�sj���Q��+��xS��-����E�c�k�u-��mxtR|�2�M�>���r��GY�~���9�F�����#2I�լ��ɍ���v��p�$�8��6δf.7dh��9`k��9z���(�慚��$.��X,�O�r�pe�2���k���.����~ǉɑD�`ؒ,��/sR5'��g�l/܎���2vɄ�5��t�r�\@X���E�p.x8�H��S�0J��O�J��;�f���A �F��ڨRAp	%���ӗ�I�-�ߎ�|��?���b���`��s	 ���#�Aw��]�T!�V�� <����>�ee	�x1��x&�ģ��9����`�o.]�Jm�����&����M�ڌ&]]/�z��B��s���8�2���� ���O�Tf��s)z�E�`M�~j2��(����dr!�+w����ӳ?]���G�
�S��L;J�]L��cTE�ԑ�A�LmҳiU�~������!����S$�U<p!i��N$���
�ŎV^��/��rw��EnǈM�ؤ,FI��5�(I�KJ�93�(�~.9�l+���Tw�7L�̓R�h-|@Vg�O:ݗ�%�C��k%N0�eTSa�/JB��Pn���<c�yRF��Oy��Ed7r`i�F�MS�.��DYIϋ��r��:Řu^�4_�yU?ތ�F��H rd�G��ǚS�C���!���^2c65*��i�f<�m�8�sVe�f�,���x��`�7��Hed�M����(�j���6�wqBj$��s�s���1F�#��ى��b�gR����w����Q2{ǁВ5)9�Qd�M��U���N\�<te��ݳ�T��^mn\���Ԭ�<7PG�Xو�#b�?9qort�[Ԇƛq%��U�q$��t-i�U�@#A�R�5#~���+p����G�����L�A�v��Ev�&#�#�ۍ�`8U�"�-7Rf�W'�j�[��6W�d"��ew��H�p��#�)g�1�LCF��d����QapKՈ2H ��*���4zR��Yz��C<�H�I�P��@;!�z��K��:#�8�7�i	�0�q.�Ƴ�v>=Z����$h㗋*s����r���AT�5q�	F�-4�LVc�3#\��uMq�b��2��b��V�
��"7̉��#	B%��C⣫���B���M���:B^�9]� �G�n4�?z�](�pK����4dޚ|0�1���E�Y�`�4:��!QOi��ǹ|�4�����T����J-;g��G�+ZK� ]�p���2��?�a�[�='Х]5�g8q�,}�����qs4��c�L�2 h�	-g#%�I�T��[�Rv�V(uC��7)<]AH�CSc��������K���q!P\�j�/�w���L#7�`���ˬ�c5e9+&��v�,�D����2f�\�`��S��#cj3Y�iԀ���D��g������~b�+ČJz<���(08pgt9�Q/9jc�<d;��`�x8F�GM&�tf���c�Z�{҈[�su�Kj��c������W:"Y��y���FJ�ǉ��$Ѹ����"��k�%����y�+E��T fEq=�!	��-hN�2�X<�������8�h����>ĕa��7�Z�6p����y%�i����+a��0�b�K�["U�0�
}���/�/,����U�O9'�9�ՠ4G���g`__z�U<�FC�d��.K�'�?��,'�'&|�@�7_��E���(��4y:V&�)m����*+K�b9�mK�F�>h~d#ڮ[����Ԅ�y;0n�K4
TN��� 0�`[(]�^9������:�Ѥó+_�CW� ٥�����Q|��[�&f����W(�Ң$�$hRBȑؚ��F�)���pRY�ש�b�uA�z��3��ZWji���ُl��h��'�����|A�v�*��٬%��d�zlީ�<<(^^]��R����:0O�Ψ-���U�b�&��e<MҀى˄�a0³�d���k�0-<�J�.��$3F��;F� ᏑZ���퓓$����a[���Bࢶ���v��hI����B� E �0%�r��84���Y�5� Q�=6����W���Ų�&N}�b}�Zf�N����:��	pR}dB�+��7�L��I���Y|Mu`|�����Ջ��$#Pn��}��#�F��fN�)Y�Mp�};���4�kC�/â2Ƣ������,Һ�'�\�,�C�vs"d�0�a-�@�U(yx,eri8�zD�L��@h���� .�%񋀙�Mi��;$��;��E+��9X�:�_6�K X��6���/|��=�X��J���r���&V	���4���3���^i�I+	�D�FA��X#Q$q�k� ��G���v���_ �酘!���G��ܤ�5?dA�>�3�a�\���8h�2� :d�F�mAiqi�[*d��G�������JGo���L��Xace���*���GW].3�������y��sf�qO"�T.����r�)wD�!��q!�Z-esܺV���Xy�C�2�
@�FX�gB�%��F����z@���M8�>6�vO�:a�Y�5����Qj���6����k���$Wǝ�lI	�.�
�a ��νǭ�	�2�#|H��5T�'D�f�B����6�k	�F�{X7SWc��ѩ��lr1
�;"-�Ɖ�z#���c���`T���sSEl��d���x�Q� *��\�@8Y�ɡ��tZ�����4]�f`���`��T(jTTh�0ʇ�s3�yk���+���v��R*�|YPIw��Q��t-Ԍ��>c��"u� E
��$�#�87d�f@�	uLQb@�ec5x�#�;X�χ8��h��2��\D��d���J|�qR�-�>3\���0�&��-j���x��Y'��Wc�G ����!���7)�X���Z3�ǦR��0���d|�R��w��g�/W�~��e��+B-I�H�:`,�i�HH�V�Bz(����F<t���'�G^�Pz0�>�t���c�p��P�>��pA�,�z��=r/��֪�\g�gT%��RSH��o7؜��n�i	�hc�p;�@F΢y 3f�(����hBi��"tź8�s��ɏ8��9cCф4ж�\ih�a<�NeF�v�ڑ�W:��C��Ԅ2O�TX��iD�@6��5�hD�I�t�pXT�s]˧�˹�˕b=OUX��8�����Gq��ʸ�Z|�l��'����j�}����g�G��1yL$��$�{�	LMk�쭫��\f���!�2�H�[]K�ŉЀ�)��ip��9k7����p��%��	c����Ң�-�#bg�0 ����A�J���ȏԶT���b�])�P�%Ϣ��Ed���e�mW!I��\�oIoB\�H�� �6G�.b�QǛV�W7WWu3/b������>%����I��C�0������.N��B��:NE��t�]�z7Vk��\n<�${7�j��K읳��z�!B`�cP��J����4=E���/2yP#A��r(�A�ؔ�%�Xtv�~߄�(���~ƭD���!��N�Ȇ
es,�NtsTq��"�Ӫ�U7 !��*���Q���@Nj�����D�2�g׶y|��^z�o���%�b���|(�@د�2C�����N�p�!��(����pd@������aR��=U�Ӎr�ʒ�H�s~�` ���Ь�����T:���	�>�E?�1?���!�{�3fʝU��h*4UȈF�7�r��X.u��ݝ�@7E"4�j��>q�����s}V*8���������p�Ojز�>��B�2Yڢ�U�@�%���!�R��z鄒"�1͡��*��ԯi���*Ѩ��v/T2�{��r���$v��F�~�Z,�{z�΋\�7 �/�>�<7�V��ѽ�kt\�x����g�\�ua�ᅥ�����_Y�B��c�,��s��~#�94E��!�4���C��/J�Fe��Y5^�Pˏ��a�"���W(M��a�� #@ܿ�nJFl��_��¤9
� (�Ē~�#�-�1��E�M�\.�����Ψ�)��E�����M������vZɇ7..o�
�)��CV(AE�;*'o4<dQ}�Z;ϼ
ͪx�j�����+O�]���.���mQ��ː�5�CC]����=�c��T�,X���p��4]�T��?
�PQ�Ś�d���,3]-�F�v��$d��q8 ����bq �?�k�T����(�.�)�#������ۂ#mMU�!�lJ�K�0/�W#�W�h�Ȫ�a!3}�څ�..g&�p�חq�����,����������d#���g�̡ۮ��o_l�syٛ�l��a��ZꞴ,8�s;H:ڸ1$����yv�ָӪ=��\��=���M�8q��h��͘ڬ��Ed���v�:�91�hEu)Ȭ�V��{=��`͈�� #6��� e�� ��)6-)X�Q�D*�:��PZ'
��0�C�E�%  @ IDATN�So���z��K��T:������&q�l@���3>�b8)��d'}���4�k!N��;��V_� �|NE���l��
�[˄�z�⽽{����b��e=%�VD�A�&l�AZ�	x"�F�ʄ��q<Y�x ��0.��"ti���$��]|����;��h�-�Ѡ�*�t,{Q>M �Uq��8�����u�����g6�X̶;=�mx����������j���3�XB�üB�K���R����z�B8(LZ�y�7?��[+ٰ�4=i5*e�?&D�d�#��C8���}r?�)i��	�o�.�\%��+��	�pN��-���|Av(��^�����l:B�l��j�Yok��������
T7���r�d���= �ԐM�QÊ��B��� �Zx[�3T�C��	kF�����"9�)-K�QA�KHV2���Ym3�����"�!"ʼ~��lG�P�ȉ��Щ�7�5n����.���$D�E��j&@pB�`�����%�E/�ͺ��������+��Г#����PS�1|��G�w�޸��	d����j���J����+K�� ��u�ɠ�/,M{R�#<k�5`Gclwl1��&/��M���~OU IM��g~���<����Ŕ?I�q�4l-�۴�����i�2��"�����lM�&쌒�u�� ���L31P#��%:�,^���!�A�9�MN��lR��8ә�Y�����o��z5��[�.���x���W�ﱸS6�?����ZԱ$2G���?���Ӗ�ovZ;�f�n77���_m��Ijv�[�2����ն�\h�$�)s*�i���J�����^�蕀�{����!()=�(�ޠU����p<�\=�
�r
j6�p�1M{6�GN�cov��k�p���������cb�k:7�$�����;`e2��R��l���Z��͕��j��`6�@iP[�G�c8��Q'3����<��-2~:�j�� 16����'756J�_�seggg���څza��պX�U#���0 �����*�hEG��E��t4$�Ğ����s?�RE��Cjн!Aj�lL� �E��r��iqv,�
�$es�~�q�����y_a
V� /^���d��U-d���j0,	��,v�]|�by�p<�[O-G���U����W¾7��Bj�^�nhN���@z��2�V9�25��xsq����B�;����SN��Nΐ���"��C�8I�˫?����X����6�!P��5r=�a�=�KK���&��8�昝���e�THK�2����o���fo�����SŊ7@�ܑ��:&��*� ���-R�$� Vz�T�?	�*[�N�ޔ����"P�%}������$P�CG1GTD�;c���b�<�$k���ݨ�~����y�Rz�7�?�nFi#֩O	�?�����;��y���,��9�)�}xcs�?|��{��_�Շ�Eܴc� �u������W.�_�v��1�&K�-}��(�֖M����p������幏��Ѵ@n�U���M���c�L:8~ih�Dr��q�����LK0J�;�&�ҢT圮b�[*�4�;$����bi3���tѺ��gv�'C��Z��\x��&��=��;}���Q$]��k����$��@	2jf˞����V�%��.8��(�l_\���w����N;H��^��*�^���^�����>,CW�h �8�|Qby��`S\�J%	�,�����׏?Y*��8���냖��H��0e.�ڥ��� ��В�iᬺ��3H�Bo&�o�\_`�K�R���B��A���� `Ol���}�F��(����i�w�7~v��f%�~����%fӰ�*�t�!z;y�3 ��b��;T Z±�F�7�!���QM�Di�U�,��7�s�E��g�ֵb��~���?}���j��
V�BK���E��e�Ί*�ݡ�
�"���&)��{�&V�`���E���G^D�_��I�����4�f��+� �e�m(X���!���Ҍ��,A(
�<^�5�L�9ln Jf�YR��#���K-M1Is�A
���+�����]}Ր��G���<K[�_����o-�S^*N��P��dKiv+6a�<cf��Gұ���:�qX5¢��3
g �3ʉچ��mມ*�:{:,���xP��Ԋ��[���0PEpK��d4�uژ��)Q{<�@��'G��u,�u�������@@~b�udk�4δ�=_�M�%c����Lk*U�)b5J��d�M(���4h�n�I䊆��V����S���d��<J������埿}���Ҽ�"����ġ���*Qա��z�����L�Huv6!j�82��Ad%��x��R���W����ǟ���BC���3�;�"��4"�4=�3\k�Dr�"$i�܈f��q�V1n��70�$;*?�@E+4(�K���	y�g�J0������������bZ-aLo�橴�=��}�v�i�Ő��j�}�Z�7?���͚�� I[!*N����i����qv=8���������x_�-NѮ
ttj-W�HF���lد+^��B�?�����ʦ˳l����?���r2M4�0�!�����	@�)h?������*��PB1
	�?�4��T%���V��	KxPl|�a�d͂#�p+=���� �)pņ(8`j0r��,MU�
�Nn:N��ٰ�֒���>��v�Qȶ��y�]N&*0abŃ�!m�,ع:T��p8�Q�/R:�j�?&p�5�*ނ�?���1��-�!��k��/o\���<z����r��Jy8CKľ|&2S�L���' 5_`Z���L_����p�pEYh|uI���;�C|�jj<&ߧ\�B2�y��q� Mzc��f��Ք�U"d�l�=�Y�s���I�yU����ޘ�$��r�!]jZ`�{6��[��l�:������k�\/7����L��4�0:J� k���"�J�j���'�G��;H|�ѹ����O�R��
�fG*K�����괊�s\�̆^�?|x�@��:�I��WbZ��"Q��$�k 	�hv3ܑ�԰�h$,E�1m�&ʥM+�.M�$,;8Z�qb�B�:�6(���z��D�Ɣ�z�,>��i��\B�ϞΌ�V�� q�|`w���p�*�����W���÷�^����ǘ����
%�qpf���C�n�B������?P�=^�,�#�Jp�����P ���*?̾04e8	�������M���p����d;��e&���d�S��.����)�����P%�T�Ē�hD��F������kEũ�ƴpqљup4m�ָ�P�g��=:w��@�I��$��ԝ|nk��%�9#�掘Rf�v#;�ua壷��ܨlx��h�VwEf�4�.%49g4)gH�D�h
Hɾ�@rT�II�:�N����N�O��+�*7��tv'�6�6Ń]���^�{�����w��������̛������$ �l0r��/��t���c	�Ez���d�`�%H[5'�)�K�fg.��⠆ə��L<���ۑ�e8p����e9@id,��N6�$/>�ŅI����YЖ�t2��K����?�y�4댞�[jx�7��NV��hw&g"�+��}�+�����2��@�q��tq\TV5�u�)�/�����܂�oҙ5Z�tN��z��a	�Zs9@��Z}���hg9����.d���_�|��C�ef�R�XIY�: 7^p�m���b#Rlj����D�}4�@��n�C�FS��"\�l�U
��=[�I�lO�4�)�)r M%3��$���x0W��
�bٰ�3,���y�iv���;���/��p�q�Пtؚ�d#$J�~/��)��ǅ<�x�!�Ïӛ���z����m���hmr��%W�?�5�[:�� ;����UB��,PG���B�k��������'�!��x��r�������tC�uM��e��NK�?1�ޭ��:���	8$;�FZ%mpi��ǃ�F�3���Ķ�!ɘ��Mz�$�}-�mHJ�h	4�N�Q�dJ�^�bQV*�zɢ7>�{}���o��퍷֊�poޟTfc�7�2�B�t���IpЀ�+�Y�JBi��������ωpr����AV�Q�Q��`䗲|p�ʦ���ËK����z�w���L'���)����Ѿgٜ	D�xu{YqK�E?f,N=k,O�n����	5�̳L:$�4;ta�I�x�^�S�%�F�
"&R}Yi�׻P#�`�����J93:�q�����o����޹�V��N}+Oኰ��a�2�k"7B,�!Ve&O��~�jܿ<��#��@�?�ȕȘj)�.�8�Y����T�дɤRj�Oi�՚�c��7k��{�z��N뫝�a?�@��R�B{�,�8�8.v��n2;�ÅQ�(i�B� ъ��K�<C%��(���X�`�U�b!(��
��1�(l-�+�~�oUf�ja�?���n��.׳��l�밫
�ܙv��u "�#+=��.��.ް�o�p6 [��rd����	�!<���ʡ���h;���:R\�"��~%śι�ͱ8��*�5�aN�t����?~t��vs�n����O��:d�N�P[�㸟�T͋l�1P�/F��k&�|R&H��̧ن�r� �Pn��d	��ğR�D��fAe�wG&Uk���p���W�.o��obn�(��s0����,[Ӊ�F�kYFmB��C�2+��]�s�?{��Wr�{§��$ ��wE�W��2}o�<��;3��w�W��Y��oӳFW�2-�T�*z:�$������ؙ��L$�`ɔ��@�8;vD���G��\�M����jS�u3���dd�g{�tKȧ5���_
�"Db")B酉Lk�kU��H�1�A�H3o�m��&��j�O���LO.�C+��2{���)3Q60��rj��g$�
�M S�2�)@��&y��T�\Io,ǀ�ɴ�������]�(2����l��j��-p�P�;Gۏ�ו'V���^: I�Y"�J�d��DjҦ�wr��Ic���Ӧ�����m��6�r�A���ǜ�}��b�L������G���� 3���49�-�/R�G����>����ū��Ǝ:o]󡎦*��Jj4�<���II��C�Rz%�K�Lrq�'q�L
�3VˁS8I��@uJD��6`w�,�n�<�~�*��mu���+�]��-�JDg�P��4x�=�0f�VY���4h�!"3��]1��6�4j�z�`��b&�&��͛��g	�vAF�V��$H�tK��@�xTG(��U��IFL�g�6�Y�$��p��\U|���;X�c�6���.t6�^L�L���g��d:�!��y
�`���{؂W3��DR!ڎ��\yu�䢥(,Q�ȕQ����JnZ{BJ����l�{A	}}�>�(�%z\�����?���ʮ4y�}\-Skp�Д��3̨o��͖R5�6�#��uɿ�|��o�oI��:�\�k�����L�E����![��F�rߑ�`(�MZ�#��Q0�%�삕�D.?���2g�� $`���M�T5��sɷQ�TU�u���)0_���熸�4�땙�j�u�,���p�&�W3 ���V͚=n"R'�!�9�#	���!ܦc�&����\5�'��T�q�z��/~f�mu�������T�v�c��c N�h\e&Y�r���-#��.�l+0�W�&��Λ�ؖ��<0oM�Eڐ��1��<W���粷����mLI�mC�[/���eܔ��Yv�v��@�ʈ�(�D�"��r�P�V�<��u>MC�N��^[=����>��;6��.�$�ѕ�Zu��O�bF�����toTz 5�����������Q*� *f
&2P�ΡK��}Z%��Oe+���� �(}+��5���p��p}M��_v�#�r{�4dF>�-*\��X���0�k���ټ���#�q�4�l(�g1�7�y �\<�h��i@���ck����_�L�(���Ah��^���^WgE��U��	\9�1�Y�,�R#3��D*g3���V+\�l�ړ��73�F��v�󸒬�����5V�+�Lk�m�|KJ�T�VV0��(�l
�uut5�uj�*���>��Ur�#Smx�S:WZEU��8j�k���~�����������͜���-�l���G,�
��൩�X� R�9��]h����7���o���N��,���}�
Oy���i��p���3���xf�3��h$��fZSG���1:З�{��%�#�~�P��m5�qWY�����o�5�׵�45�}���{�վ��:7�/�W�!I����Ra�bKr�ARh�2�!fS��a+�
���� #�3��ng��n�9�FsIoE��E�ɬ���4���z[�
D�ks�%�<��$HX�'��;�(k�d�)��D���hw���2�y+]���zU��%}�)�V�]��hb)����N�6Pk�4���BV����jU��������d�vee��[�i	�����-|z���a�es���Ɨ�k�8:�C{�U�\k �%������{�tֶ5:\�OK�j.#1��'�6�Az�d�J�*zȡ�L�TZ��rW���<9�K1����9�[�[�ҽ[�6_�*�!����8�.j���:hʬ6&�m����h6ɮ" f��Jtl�6���E������u�U�ʲ��
7��Q�jYf�e��\��w<��婢���˩�2R.(��������HTM�r��h^6[�<����)K<�-�`A��U�[�E=�ʙS����*����$�M(P��L)X�e�`F*�N���ur�CB�W�r�7�T��f[�ѿf��Q0���&��J՝�8�s2�k��e͛���Nr&�9�u��b����4bن���lD�lC���5��Px�yvl=�X���tsH��`[:t(��:d��C�Q9�q�>��b�4���):�hR���V�[�;��l6��9�/�A�&��a�!b��N<M;P����R��G,q�2�ML�2S/Y���y%���Z��aIU�
�B\K*M�lB�F�,� er.�#��ȑ9����. J����h�ij I4�sHL�'��=o��_�_�P�4�9�%�/|�dPF�ڼlmT�x{P�=|Tsx�#2Ֆ�T�"/�l	/�����SQ��9��Bc<��kr�1#����C([�l&	//r�H��"���K��������8��X[��$)�4?��@�o��$|��d6Z	��F+�M'����q���%S�|s�r5�=��\��J���q�O]6�����[M'��l2RU���U��.[Mb� �T�	u���<[a���mmu�}�uH]U����F:�s3ِ��V�Qa��zoy6�I�0[�E��|��˼I��\���g��ѫ��A,�Y)/Oy]LD|���}�ٍ���
��cod�׹�!�X��Vdc���dt���/�D�*S�e��MWU�j�3�Y��_u�����|[3g��8h����o$�I5Ъ(���1�J+���0`�b��`΅m��mh2�P�nI]B�0��P{j��ZB:�*w�R�h�X<YWWhl�ñH���3��c��j�<�vU񵵥�`m-_���-�٣�2�]�R橩����4���}LůfcD����\����0����5|���+�PWW;�d2��v*�G$b�զ�&��Lė����d~6�
�---�������%�7LLδ4�Ը��K��ɢ9��Y_Z#�|�a5a����
�07�ծ���������LPch�7��ڪ�����:`Z+sUe#�Y����Ĭ���j����(Ue3���ن�@CS�Rh�]���W+���[�.W���`0�������D��0$�����=k�R:H٪��@ft$3@|�X�d�;Z�V ��AV��3��k�|ϛ�҉xlbb����B�e���E��)�d,�M>\_�������H4 �HGg� �f��gffO�8�7%�K�s󍍍]���N����>}��㙝������O}������i�?޿8?���+���\�>�0?��yCC��ĉ���������\"�?���?s�L8#~�e���٠��?z�h4GVV������<{����lod��ŉ����q�����T6S�wy�|���Ç�]j�����c�����7Μ=u�̹�����@ p�x*��q�Fgg���b��7__���g/����O����W"��?���\Xt��E�ɱi���gS�ăG����~X�����cz�P�|�7Ly�޻1��\0jm}��2�����SEd�\.��&��ٱ���mKS��G9{499v��͋�����yu���#�����?x���Ç{{{?��S�����jnn��O~^ߺy���}�ч|@��7� �:k��7��?����c�psװ�*�П=~���x����C�~������;���_��_g=���n߹}���}��[�����Ǐ>��������_��?��n�/����_��;��i��~��K/�?2>z��ݞ�c-�d���t�}�ṯ����gW�����������L6|���٩�3�������/�%>�^N/�%M7��j��������S'OE=3��#�6�+#K���?y�����y���?����>�\�ܽ��XO�\�n|��o	7LNOݿ}��;�4Rb����o5t����
������+ì�)�Y8c
U�roZzW��t<��ѭ���L2XS����?�?#�6�K�˃���O=;����g_>�^�l���'�
-�<��\��>r=��9P�J��:;������ۘN=op��U��?��ލ/�e�@����{�����=�ٱǰ�n��nZ�|t��v��z~���u��t�'G޻��z��c�3��n���&�B�/�}YS=u�585x���e���*c�CwƆ�u�U��L��^���ջ�G�|r���vwyb��ՙ���5w�zƟ�<���S����n���l�n�g_�����]:~��cx����@SmՇWN/L����_w��������G�[5��n��n_�Cs}����V��<�V�^��z#������ɣm������ek��}x���V��md��P� ������ԑL;�a�)Y�A_#�Q�|��^w{Õ˧kk+�>��;��������ܺp���ю���z��^ow����T���9u�����;���z-~����Ƚ�_�'9�{izx���F_��_��n�����C���Wm��珕e#�Z*L�4�Wݼ�E,�����)�~x�;��ѻM��n_M��?��g�G����fqv��9~�c�������W8:�6�����ąS}��~5�xd��#��~�F"26����w��+4=>�r����F�g_��V��w����ԃ�_���ϝ�	�O���&��G2�ು��ʲ�>z���Ƿ+�b�O���FG�? 7'�:j]믆�Wf�����Ã�f�f>z�l��>�������GV����_�t�8�rt��ᮖ#ݭk�hb����7?[Vr��>��A���ٙ������hY�W���b�1jǏu��ռ|1��壺��?8]��}틞����+ˮ<~p��_��Ǘ����~�\W��O�uWd����{��\8�T[���5�u�{�\w[��𣊵�{�O��ܿ�eh~��I�P��������<C���M�?�����ὥ��c��}=G�F�WBK'���}�bp~v�hߑC]��S�;[k/�9�095�p������+�N�z��K߿|%�߹�My&���ȷ�&���^]?{�Dm�{����|���]�����.\�w/�ˑ�)�᧏�j��s'�7>���0���gX!x��Nti���g:���#�gFA$ٜ.��t�v5O?�q��s�̱Xh���oz:�?��R6~��8֝�_=hn�=���^=��,�,�B��d.G6��mfQw�} �j�����lmL�2���+�s�����2j�c�N����9thiaqn6��D��a`�I2�:��o>��~1w�䙖��C��GN�<�s��ȫW<=��{��������d[sKC}-�����6��˗�S�����"8^��ܾ��|��ի׹h�K�X����;s�b޽���5N=�]�ׯݎF���\�x���/��c=G�57�߽�pq!|�����'O���;��t:27;���Ӛj7����6��U���<����ݻ>w�;�,͆��)�Dol|b�9���N>�9::�	�ޣ�W���`����h��$���G*k���S����S��ֻC/�������adlrn!���_[��?~������<}���frfnfv�������r�ٳ!>UF��< آ'&Z��*��F�8:}X�Y�O��v�ʐX�]�/f�R"��ϐ�����QT';?~���w����������־�ޏb��[7���v�:�AY����$̞޳����55�S��p�����X��+����s�ٳg��/|P^U����G������/��==�={�}��������˗?mk�{�t�����3�����^�����ˇ����^y�l���K�]ǂ��v�}ǈ:��?~�4���~4���/����~���T�7_|�m�����%��|�������?�p���_���>�Ql�����|(���̚����zͧ��lm����������SS{߃'#O��?��?7t������;���Љ˃�KWｸ��*����|�١W���pl>~���ѳ�}ͽK����z`������O�eG'n�?�K���>�������H�jx$���DUu�|�`K�K{52��� (�Q^�ڹ���H�.���4�,��~|A�{ ������J����3�K������^�b����s4�>00�����s���d<8�x���O�6���.`�>�_��/şO}��Ǖ�uφ�^����-5��p$s�����ǹ!���W3KMͭ��s����74�WxGF�&'��������׮?`�>����?~�����{�,��έ�'�\�յ�}0\�=v��o�z���ZMK��Ʀ��٥h��6БH�O�/,'�;{7*��#��Zk���J��S_|s���PS{��t���X,�~}/����r5���S�+d'��Jd�#񲛷���й�S+_�x<��X��C�������$@MT&��+Ѳ?s?���?����qgh)��Y��.��>x���ݨ��
=�Y��U�8O,%"�"�_&���4u;KoWn@�Z<T���?ߖؔ�Pى)x)`q`��d�J�]X��#�!,�p�=��$W#+�g�1%�p�q4���J��O�>���w��V?\����4���Ï���O��?9:==�8<�]�x��E{G�R(����Rh���Og�^�M�/���0�ʼ|567�5q.n�y92
��_���=��	&�Y�
>9=74<�����������x,��'3w�E��_����������Bhdd|fv!��LM�=|�ly9�J�NO�ݸy7���MM͎O�ONr�utzfa|rLC+��c�ӡp�W[G�o߾�H��dq1�(�!�K��D��՛,�.æu{.s�7*�{�a(�F���O�ɦ��
n�����9537:6���4�S��%g���Fh)�#�N��:]YŎ����3Ef֣r���{��	>�a}���2�'�o c��!�Ʉ���H�Y�a̛+�@���ܣe�R��@l6��+�������?��C"a��%�?�(PQ�����ss�Ln��^ROZ���y�G��Е��?
1���a$�=8$�vB�=~/�����Xjdf~~����	3������:���X�io���=mycc���r���,srl��f!F�R%��bsqG�߿��L���!߮�Һ1�����d�,H�<�-�m=	fZ�����Φ�h4JR	N噚�fڙ�-|L���'%���U>�X[�'/^�'O�\5��0iL����-���)��0dI���;�
����9�@=�����c������_���A���:� )l��SؚZ}ĭ�,c����
��,{��+W����P{��%0,lܻu� .��y��"�h���ţ�?p�|\�O~�rSϊ5��i����6�4���� I&c@������$!X9j�n�
���d�W��s$M����b���'0Yc�Ŗ��Dkmc�'[�j��W�ut6g�*y�!a�(�xPv�GW��h�m�E��T����H����j?�uuݳL����#�����y8��p�>�Z�j4��m�����H,��r�>�k��8�OKˉꚆu��Vm���P������Nd��J:��H�m��_�N����Ro*��HT���PmXi���^�G.W���5�e�J.e�g��C+_UQån��I3�h��I�8Q��� ���lFE�H+���´���6������g�Ⱥ���YM�k}�Q�m9�u�	�A��� ��H�V��d�Z<�2k�n��a�<�^CCY[��k��z���>���oh�%O��s�5��3��BB}S������j���e�p�����w�CI��JO�:����2��/�㥃��-,,P�[[-/�S٪d��\�XW�vo����P0ȵv��M�ՙUV��hl�|n��r_��&do6\�Z�c,��&>���R�DM�������`p���o{��� S--́_2����r�sr��̝�3=Ů��h|�d�qǲ!���k"�
F�K�j���6 ׷��R��Z��4�Ț}( LZ������-����Z���b�z��SV�rT�g*+��T��yX�f�I�G)h/jj�[덢�#:r>��8F�^-��ϣ�Z�̰���E6��4�^���g?�>u��l������l���}ω3��觭��l����!.��z��v{j!̇G\5��P�����P8����2��x����b�!03�H����Ϫ,��.��4��<�·Y���\0�z<,�V�qW_u������(@�I��^����kј|�O�ָ��Xh����t��L&�6�ֶ��O���;'SP��X�>P+{��X)*��6ʢ��x�8>�J%c�px����&�NF�s���=�J���)���OjJ�@�� 2���4����[��`C(�Y}}=͍��d��CGSs4�*�pU��A���:=H���f*�w�����>�A������;��z�!4sv�9'���]��ϡ�u.�;t�H���&�Ƿ����4�\�E�n����O�f�h'*=#j��H��YJ����`��F�� ����\������n�i�9��o�^X
����@��FSK3E����R{�/7��3@��u�D|�vd��X��q[,���>e��M��5.7��n)�?���qO����N�Gva4�42'���N��(�TzCD�LgQ��՜����%�#�o=�����pf0F��I&3��l�(Y�>c����Tdt}OώQö��h �D�`���zI�̖��*�+�&���\�Z�KF�t�~�!F�T�(���8[a[��à�e�W��<�-�0�˟����z����g�*�aK���z��2z��&��{�H<�{��j�0��E�����/Ì]� &��O�]Y�vW�{Cc�����Oh)b�������\QS����+�:�]��$e��.�U8njl��� ���� ettd�����0�|�y��^6�) �J���+���8y����ƍk�鴷�fa~�����,]�����'�9�=��u��w�w}-������-r����裻Pg��G_�X �)��\��h2�$hۥ�ف�qw�=�v��W(����_."��N���2~�{���$�rғS�:ű��9X�WXDDً-̑M �q�H�I�o�]bl��c����b�g��/������;~����PWwKKՌ����/^�zu��-6&���1�J6��!�����������O?�����>}���u���w�\���e<��C�������ݾu�����lgl����/_���0�1�D|&s����s���p(82:�	�ʦ�t2wzYI{ SL"-��dDe��t.��h�,/bs8?W��:�QC˲���-�"̮{-큂�Ts�������Q�-�פ��E����L)t,�?[6/�ڦ�[#�Ǡ�M��5�r(YB�Qb\��iWS҇�$x�vd�Nq޽nl�HG�ҥK�~�I��>�)|8)��������x[[������wΞ=ǲ�>�L������?�	�̘Y�x��g�}v��%�M����1�����}�G���֭��������? ���ɕ��]G{����WV�'T��0��+�� "�D�f5��L�ACD���UīFn7˭q�X�aْ/"�Ǖ��&�x� +J��΀���+�
����*Q�4r�$H3k��j��s��@���j���#/���hh`�8ZBLu�Y@�d��%��,{���}TIB]�Đ*0�P_����a�~h蹿����Qi4������.??���O>��v�i<��,S�t�V�i����9��7=3�l�t3h�W��	d���%�	��
%dJ�,w)d��J45�D�@I~�̤��{3�(��y��]���:i*Lp�ZK?'C'݁��	^gSo�Hx��(oT?s}�Jo��������	?@�?�%�Wx\\�&>t��E�arJ��qJY�'Ϥ�nህ>(�ޞ�E�#�h��D zl����t�[K
�`/���T<eZ8�f�ҭm�~�ᑾ�3ӓSSk��OR��L�L���r|b�H_o�ɓt�o�_�y��3�DY��x�������ºz�.�th��i0�-�M��� cG�����&HA�d���D�=f�+�3�i���&���5r��{��RR�d1?�|4Ov��-����@0֗�#ZM�̊����ðos���P��#�3"l���q|��ѣG��&x��4O֥xL)��`GG;�7�8ʋgv5�����Ç<2#�Dݸ�:/�X�w��4�=�a���a*������ǏG�/��,�X�<�ݹ�f~�
�c��Ц�*>��"�S�����dօ�T!�;�J��t3��R)5��U���Ͽݦ�ɿz��N�#X1�CF^���/��y*�Y��ڌb�����:r|d2'';�ZC��oi��v���	�fWO__�9	"���E.,bN�i[|���{:�:��hk"�l����BKK�������*7s(��z5�t-HBmPҀ�ѣGK�`cc-#`զ��q3�
Fjı���z�2C�_:��,�p��W�t���;*�\$���Ch~Mۢý�[]�!���r��0�eR"淕zO��uh�AE�߾!a�cx����Q�l+0=��x�+��9Kr����&x���P/����'(a��d ;Y�a6xҺ��U�z�Ae�%�*�䅢E'�`�0%e���X��~�����)7Y���$�J�.���#=?<�7�� %dy��/^��΁]�W�9[�L� UQ��
� b��F�剜/�]��[a��u�!�jPŅD��B�꿥̃Z��lƐ��@?��'C*�DA*�/�Z���Ƹ�*c+��3: @��F�?�^f��Q����7&C�+��3N�G����l(#k�P�ȑ���F$ 
%��/�3����@��]����R�99���Y^��f}��+b���@5	���j���8�~��.k�K���{���_���L&���*�7���l��`���-v�����7n^�M{K{S�)�7�5�?D�6�e�J��8�A���/'Ռ�����t.�w��$8����|�m*�2g�m��;��ISdN�}�u��V5� ���j�$��:�SI�F��L�.����%�(*�T�=Dnj�H%$���_ D�u�-��2`����F�Q�#�=��@=���NniF4�b>�`��w�D�fT(���=�~�v��1<<<�h`ff:O�b�8�%}�1��5�P����/�z�od�j�+�6��k&�H�T�X<Y��iP�lv��L�VM	K?��Ћ���c  @ IDAT��>�-�t���K�P���@Ҙ���(ogd��-`�H�3�,�HagWgfg�(�<��sy�敔d��7�i3g�iI�1Y�E3���$���1��.Hڨ`�[��	f	KF�(9�-`��G* �JUf�qa[����1	zM�Gq)�@od6�����d+>�hr�[l�i�,��d�neb���e���b7��� �>�Rt���w��'Z�?��񣑑Qf�B�A��-�H��k~a�I
��3����,9ޢvvn������(N��l�R���T�\����d��P��B2�me8b*IA"wxD�$l��T)a�C���j��w�i@���b�Q���ɞQ0 N�ی$m��γ?���CY1�on�Enb��?��LO�뛘��7�!"�#�fg��¡�<�3��|h�<~����fjj��<>>���e/��|�~�2�%����#��
}FfC�F�8:M�ѣ���9r��I� X���d��;ArüD��h}⢒�e�	�aɈHN~��F���x��p�PƏ�&(P�d!"�%�yãv����]MF��a�&?����-Q��0��"D}���%nD	���--��5��%͍�= e؈*H�F�@4 �sr������O9�}��eIse������(�	ZX���C sZ:M���<PO$F�QQ����p3��	z�]��
| s&I�Шy�����
�M��5MdA���/���j2 6�A�_SNB�L UL�!�h��!4��ƨ��Lt�p)i&Hi�r1�f��f]�J��`R��BR�髠1Y"�q���)z���.��5Wgg�7mưL��^^��͜����}�F�"r�x��'�5"n�J&٠!�3WYB%�̡�	���"a�a���9�ه�T)}2:�PZW�J�}���鶞86)���6B�"�Ž�Y����ˬ�J�D
W���S��Gm>�m�Nm�i-�1�X\^
+]`�����#�4Dɺ�3��Mo�G;�	���p�Z^�����B_٤::����jN �i��4�L�p�E2!|$��T�6��6�N�]��ǈ �M�B)��?v�"/�/~Tm�Z���o1�b�k4ův�aOb$����ToQ��03����	�����lN���e&Y ��i����L��c��|u�.	�~��r,&��R�������i��!hB���	8ܹ{ȄHfUot�	�#h�H�ю�bp��$�-�m7�8�g��65�;s�O�=}�E�m�/-.�꒱ı޾������R���`����y$����9si,�ޠ!��A$fpb�� K��?T��	th�@����E^���B?�8RH)���!�(�k,���d�DX�&v��}L*.��u���r̠L���@	��S��z��f�) �D�6"{�hq�+z��2�LbsOy��)���"�0��'ڒ�{�zA�Y;�x���8��VKS-ߛ�9����?��ͫ~��3K��x|2�%�����B��'���a?��cϑ�aV0A3���;:�p��d<�Hr���RQ��*D�gYf��$�@	?N�ԗ��@,oȔU���D�v(a� �ٖ"O��_�T4�C�΀�ǯ�����M����I�t�3f\�Jo�����Al@.Bˋ��Ǐ ��e�����)m��//�]���0��Pp~vz%2�𘺧�N�8=l�M'�_<���r(�uظ�JDO����+ܔNύ۠P����wV3��JNM�se?_�	'������.]8?=9�����������
pW�q�,iF���K���"�Y��Ӽ�%�4�L^(ȝ����J`[�D,bd\'�ˬ����=���ߖ�Ξ΀N�3��5���k��;11�ɑ&����ӌ�6�@A�����'�R�(��3���q���pQ�ҪE����.'���\f�r���Ų��� xDW�"O����\�'N�<|�0K�l͠��<1&e�����sӳ��C��'O�;XU��k�1�P�"W���C������־�>i�+d[���f��ٔ��X��!�e��ڍd����R� l*��3ـ[د2b�bY�!X��S4�Q����o�ao �l�K�N"��U~
��r��EO� J�e��\^�33�/]xI��v���mV�>�X�g\�G���\����Q[���
��<e�!�g<n�Rhi��0�� ����.�؁�P�1;,��޿�&�3�����x���a ����FGG�KK���/��IO?W}\�h�����+���p�N!ZFvs�淿kmmf�첞;�l�n�<Zg0m��rXm�UD�r��ĐHM�G���̜�V���w��r�I����5�r�&(���2���D�!S�F�D.F�W#��),�����8���q�BCLMM��9�b���M�����-�СF_�'��s��nk� (����Z�ߟ��FGF����jAyÊ��|@��R�����PKˡ��k��޾[f(��a3���ɩŹ��������6� ��1J���]�~nh��U6^�7�����hb2ɣ�e�W�]�%��L�&�4iD��+V+����d�78�Cf���
hN48��G�!Tz�kf3��P��k�Ms�(t�pj*�ؐ��88�K���D8�DX
�hzj�f����3A��l�)cK�8��&i4���]�n�Z�ke�eƄ-Qӑg��pB�(X��;�H������L4�L}����~�J���F�	@�=�f��~�FJ�J{��R:V �b�P��#�o�L�-O<I����@"�j
ӽ�m�m��^��@�I&�E]K�@7��2crJ�0*q�}`��@z��J�,d�J* ^���Ф߇���	Th�a�&"b:Ti�I����Fn�` �(���t��-M������<
�҃�p@��s���&��̼j9yFn*+	�[���Q6�Қ����^�q�7�d�c����4����	�N��!S�D�V�*2,*K����<�9V��Ҁ�MY�(�E+�����Kӹ-���
	ȃ���v0­�G�q�#�+GD���i�EF>�~���=P@�`(]�T�1���M��� ����0,�VS�X��rh(8����s��2�dSC=x���z���b���%�	Iq�0��"�&�qm�٦���i�d'UU���jC�N��C�3����^G:ڻ����G�٘�b���}��t�mX��#��� ME�\���h5�d~���TUS�MX�dӫ��.��כ��9��u�8��		�7������D�8X:����S��d�]�R�e!��J�i��! t�-di��	�q�Ec@ -�Y��u��P��Gq��i����a\����%|���[zC(������a>��Qi0B%Xэ2�!c1^����J�w��DͼZu놜&b���ŋ�i:������z���Kf?���#G���\ڸ���d%!������FFF�z28��8�d�u*�]8�������V>���W�^]�z�H(<M?)/ՖA@�l���"Q�f�f3Wy�1T�s�ZL�ɼŐ/��T� ш+�c5�|G��vAF��B�����,�f����M�˙;5�%��TCQ��/#��@P��A#�DE�+���p����l��̜@!��!,��1
i���B��}�ɿ���3�"���_�7p?3?�L���CY`��@ɐr���͍޹�h��{��uzb�=��oݤ}������ �5�K�H$z�ܹϾ�9�Ł�ddJ������w.U|'�TUrVW�nm�Bh����jg�K���rf��%Y�S-S�d��Қ�v��9j��O��#:�JΪ�+u�ɦ�xm�\������
�q@M[F��h`��n��G�D�1�Hc�#.5
8�!����2�,Y�b��1�� $����Ř�!Ѐ�c3>���#�;��D�	�����*��2;�<CE6��T�G�F����ϙ4A2U����d
��w��;�Ǡ�m�H@�g�O�I'�H������
}԰ru�4S�xE�I�(�
9���)qBoz�R�0��ͣM����2��(~"�ƙ �)�"7�ৃA�l0A�`E74��bZ��.(Iz��9��K��$���(�{��|�C�AL�o��D�=Qq����9������f�9/"�I��������l��裏z{{��
f�^��'C��̒�**X��G���q��i��T��}�8�zAlm����-�Bg�.��	s@�93ނ9��[Əf/�S��e��y,��b]O����H	԰�\��@T���ih����{4����6��� Q�܌Ĕ��o��t&4 )�|���8�M�b�|er�6ڑr�'�i	t�#���!��gD)6�q��J ��O�~�ˀ���d���9
|,���qR�8��ٳ ��+��3B�gB���K@
5��s,X��䩓�*f�h4ٿ�\	#V��̥1%A�JX����%���$�E2b+����E���"�\��q�Ɂ2��a�Cf�
��v�lJø��Dͅ	ƕ'|0y�1��2�Ҥ�^V�$t{Y�%���B�Ep,�����pom&���+���!�	�*��qE 
�8mmm E84�|��ȹ��9La<|��#�S����dbb���׮_'qlcdL�����[�����gg����.��D�'Ư]�v��1T�
|��rV��^��?�h�nmv
o��rɆ�.��E�
z]N�J��]��}I�b���2_C�@@�����i2m�K;�=���72�޵wu?y"�M����Xx��y�SS&�Ȟ� ��fF�������ڛL`�f����A��N���\����hni�ßFCߌ�Jp����/~�xR��X�³��I�th�)����4R�y��$��,�<|��n5S�|���ƍ�)��nݺEyӼ�&���|�@>C�-{-;�D'���������*x�A(�k��d�UYȘ.a6�����M�Q�N����7��m�K�J� ��5��� �3v��N���~d�))���SV��p04:�j�k6o�ez��f��h̘��G����	E��`�b恚-^�P��K�[��Y7��7�x�΂�<#U"o �f�\\x���o4�"@y��Wl@a�SKC�T)�Q6UºA<n}K3��H��e�VԝaI��s����S�N2k�F� �^'3�c�4����CSKt�z�7eA�z�?����4��ANLO��k�=���'}�����X�%��MΤ�7��F�ypl#\�	n�l�i�&秅!퉑�mTz�oBm�D��Qvra]��~n�\��1��͕ڸ[��p�7KCr�L`����!BcA�5�����f&)���'GV#��LaMCXQA'��pD��!�&c��$ۀ� 兩�@FR:;:��f������F�N+%G�^���g�Pt�s�����D�!Jco�k[�ٰ���:L�M�����ӷ�-����f����1;W���
�Z�
 \�8��lX	�@�C��0TGAzl��8ӨA$Q(���V�d2)-�0S��+�Qi�b���.��/[���l'�8�e@��u��e��]_��t�s�O�b�L�j�K�(N�׀�H*�輙���24&O�Y���G4�	�^qJ߶�&%�Z�d�K��]Ly�$e�!~l����%��'�Ҩ14�<���G�S��0����A }��ܞa8H�R�5p�����N֘��\Do���0Τ*������{J"]=j�1KՓ�Q�����́20���*GmJl��)��蘒��,�Z����[fg�-���oJ�@J�`A6��N�x�p�R�@�P��>m5_g*gk�b�ۆ̩f��̍)C�l�/htjkC)n�[����Y�X�=����lPgu���,k�#�*������S���p� sr٫���h+�K&T�s�.�e�Ȳ�1r�Dْn�P.���G���Q�o��+4�^�L݄M�X�P��&�[H!9X��<5�v�d��,��Eզ��#�P��7pɬ�99hv!��hL�e�a񀀤���?5Y�l�W��ͥ`���$j�:R�k�����ur.	2�z�� N+b�v�&-I
��D���� ɬg�3F�O�1�B�+Kg�L	��K$ ǧ��Mo-Y��994��6�tKR�u ZB,�2P�G4}��j)|0`e��v��D�WH�I�4~2r�� "�S��ւ��Y������%���'Z*pI��
���ȕ}5����挃��+�����].j����Q�b����!���c��#4���  b�_���6L�Sf5�Z5���*�%;|�$�\2���M�RX<�rjb�Q��n'"5'y+���,��掐+]Fht��&�Ҁ�x-+�g���/Ė���� �;�����VqoW���.<C,v�fs��#r�*�?U���ɛ�Sde�Pw�ɭ��A�8�z��*���L[�̓���^qМO��?Z�{�g������K.�n�,h�����Ըr ��9�K���N�,��#$r���Q`�`�ca}(q�����u�,�Ύ׃L�i" >Zܝ����f��Se��.�Ͽ����% zT�9E�[{�`y���(h'�bn���Xc���QdćQ�V�Y�;c��r�١C��4�f8���C�҈��YҒ2�_;���R+�-�DC�Z�,)��A�'q����J�̆����s��i1s�7��Z�z{��=qV�i�[[�ԉkg�����	D��V�;�}=�,zf�~�SG��͕��l���iR�l8�&���+��U.�2�T�V���v)>�aO���=�����S۷v�ș�b>ŒQ���fg�d1�tUv��R�����9J�Lm�$xT[�-O���~��� �XJ���a�e����%.vP�)b����� hӀŔ��z��N�8sr�����;�I15�P�NˍPN�L��J%`�I���<U�N�ı���҇l��P����vI���e��6��P^�XS�XqFSඳ��S��"`��XJ'�����@�
�W�e�1o���#�lݍ�o�ۇ�������t[ PX����*6
]AV�$�&q�{����b�<���w5F���z���g�� �0�n"��lä���²u
�I\����q�������y$�f��TH���%��&�q|�$�T=4j(&UȜ6s�1.��w�q��)
�aI��.��NF���V�$��(t,��ԐP�=����[bx�,	E(d�p�V(C���y�a�kE"�(��Lp [�Rz��%�@�4�U%�TbsR"vd�)���O�2W	;%�t�"d�բ�� N{/^k,�� Xp��XF���Ho��PVC@n5�x��؆%��GX����>��U��-��Ck����<�-�5���^|���D#��/�$�0yj񱥑G��-B�-厧�ط�(�IL�	e�T@�=�(Z8l@��G-u�t�"&R�[g�H1c��(��Zr�����A��Q�����3$�A�n�FYpJtjj��1R�t�8Ըj/z�"�C�x�A�x��xC䌍A���ҁ^�-��#���ʴd��d��0%���G��!њ<�PÈ7�1�`K��T���r�Cr58A��Qc�vͼ�Gݚgu��8�d=q��S����t���4^D������@�$�[��|A����^sD_7���.(a��C@	B7�W�!�-2���?�f{�Aa�q�E�h��G�aM�4zK����%����3(s�{�9{�!t�B^�����s��8��D�3�7�W� �D��qvf�e���X�Qu������w�_�P$��6��B�yonns���k�Xݖo��-�	�m����I�La��P|�H�����̱r��n�g�B�"&����>�*��Y�Pb �V�B��4*j�`/-Ft�hyeY�G�����t�xK����#G�455�Jv�ɝ��8��!zrN���|(P�tx��	1���V��-lؖ��e��(�j_�H�*�a��� IWN�9B�9^�*ނ!��r��!"B]�v��xyQ#yE���?���ag����p��ľ���>��,x�X������!/d�	C��0 Ak��Z".��pW>u��W�iy�J$	�?~L=� ��(^a��*�@�VP�'N�(&~=ȈIY�Pnbլ�m��V0���*��S�����8�[)Ʌ	�B|(E8�z|���^ij��'�4�;0��_Q�h)����E�'ME�C���:�;�>н&�qG;�9s�����ǀTˊ"@���EAFI)� ����UsY������!2z��(I��Ƴ �nU�5�{�+�3U�DJ�X��4����J�$��J��6=���._����y�F)��?����Q8pX��ĉ�}�$�~p�1�0�>j{�Ń�F��'��Г���E`X�#m.6آ��3$�1~q�L�>S� �����AdB�D�0���l��,�����)u�����}��d�A�P����C��Z�=en 	�!/�Z�gxR����ʖ�=��%�2kNi��V�
 (W}�aC��������2��br8��?W�Q��0s�zs����5���sC0ʝD��0@���n;*���L@�?5��n�$�d�n�ɓ'4H�F�j�Ǳ{CXkJ�H��Q�b�&�68�C������BӠ��t�7Ҡ7���^���!�fx�3lpCD�+��3�Ȕ��FE@�P�g����]LI�����-���bS����@����b�9���fJ�7�v H2at�A�-�Ǔ;D� cz���lh�Fn{���(��`<���#|P#r�9���>ˉ��U%���S��{JĶĊ!�P?C*�Kސ�f�fx۰o�I�y>o֪g��q:�@��QS���D#'N���k�$��&��������qёfr_Cip��q� ��$K`���a�7��x�ԨS}��GA�s�� ���m���g����7d���+��&1�y)��ȸB�!�K�.�SbN�R؈n�	@��jB)̹JW��1�wʜHwɿ$�4�0���Q�H��D×fP6��wk)2९�C�����A5R���0�b�fM)�N��p8��n����/�F��R`��>=$:aL��i&&&��Qk;Ƀ�� ��(���遁60G��޽ː��Y!dV���#�Q@��5v�XSd�b��`�ʷZ$`�+XQ�DG��WDZ�������f�j %=-S7���~}6��"W`Ha�!R;_7I���\M�S��6�}�LS�ҦC�>#�6q���F�WpL\Tb$�ĉE��W>���ŨT�)C�K�ol ,J�:�oh0Sp�hD�g|/5�d/�
�
����.��Ȉ��%�AP��I�j�4����t�����v��7����@Ab��l�_�U�|:��/�-d��U�x�e��g,�8��{�Bõ{��dā��i��2*�G2���2��<�a��D՚D��G���^�-��&IK�ض�{�z�D�)W����;�C�h�Sa�&:�Q���/՛Gނ3��]2�Ȕ#&ʌ��EjjH�v�^�蓢��,q�obWA���M)-�_�"���C�M^�0�>~;	F�H��}���0AL6����*\1����Q](N0�뻉�������$�U��P��P� K����֫��g74DJ��nk�x�&,4��Sv�����P���R��e��%S1a[J���H�@nmCi����>��b<�W*X� gj��'/<��W��}�X�Ĉ��-� �f��&bbj�T�gƴ�ג^A�m�m���P���QcDG,tSh���e��\�ZM�Bmg�9iJ���߶[�����#�'G̜��I�&�
���3F�Έ��e�lOO2g�LK��ׄ� ��V\i؛&S.��)6����l"#8�������a8�ӮhqD"�� +������ ���G�@��e֐-���q=:��rG�4�L)�hSE�<�2�����)Y"�D��3��t��#�G!
������<0�"(���|D�:�H���Z�j�&.� (�T��2�=����������IВ-����e���Q�9�Q׼ͨk�mJp�/F'��~7#dN�E��.g
��8|=����X��*�+�,̳��Q�VuῧX�22I��g3�� �"���S"��5{z�4�B��?�pKV^$��O���s�-�S� ��綦�A��}�W���,+<�Q�0| �c{��W�+�Λ�A�֏�;h�YZ����\$I���S�u%�Ȕ)!a������3�����Q�N�M���]ܜ}�lYC�Ш(�����_iI�䌛�̩Ig�؇�D<�S6(h3B�@`eh�P�w� *6�L�{�ro ��%J�@�Y��,<P�[����~��i����Zt��*�UK�N{�I�^y�-��ȝzE� �`���'�iL�[P�L;�>�L}�G���۞AFDC�4'(-~ZnT7�8���zIM�-5�]M0��O��w�����R�N"���S� ��͛7�
�����7�F��dW��1忏X*��p���C&�Q��궞t��'�]�M��5�D��
Dk�Z��UL�t�č'q�D*v�^3��Sɀ5"�@���b[�{r�Jម@|�|`��dN�E~q�3��x�
M�4��|���[��A8�_k�L����6��������+��d�R:hYBA@;Ƨ�	^��4�f۲ W��PN��l8�w��}휑I���[�B
�e��zZ<qS�8�+���xr�*k�̆�{u %2e������B�'�  �o�fw!��zHc��8ˈ�ԀG|A;_��T[�wó��5�mD�l��66>D���\�?��!Ҋ2�4)�e�y��:}�Tb���y��ɧ
b�HE3������TY���n��n(w�9(>�X�b!���#6rF� $������(�,8��))XQ�A�DDs�0�{&���m3ނ�� �R(�Í���}�L�/ S�?�&q�!��ψ �����Lԁ��%�����% �GWQȉ�1"%'@\�<��F�K��b��;��m� w�.E�A�� ���O'�0������ Ct�����7n܀�ZMFإ�k=`��f�X»�u�m�����}���O�L�H4'��� sT)�	I(u�[ ���n�k�^�����Y12�c(2C@�;	�heqF�bظvv(�bMa����c� �ɐkG҆��'g�����/�}>###��&=�'U�9�<
���Q3�N����	�(���ޢ5��q���y�8��!�m���2Yc�$>�	��[ʞ55������s'�@ЀB5(a(�$bb���`��CBv�Q�0�4�':�Ł ����A���A8�(������ER-�?�]d�<#�W���A�E�`��HΔpp���b�6����ڻ�6���y 5�a���]KZ��0�'A�aw���
n�Xd��#������)�4,��yKX�~�!DC��RC�')A�TD��a��k�w�5��i�o�J�[��L3��5�E&�   �!���RiiF(8�8��6e����� �c s:n@�
]ʂPj��$ɀP�����x0w0 #K$N��"b�:��X�5"M�f���ѴR�!G��<��
O�+Ȑ&	b�'�Μ���=�2��O竽�;Ör;�$��PQT~����"|^Q��Bc���)x�*4�q`��'���y�Q v�OD��Q�|��;�	��v$�4�32mqCp�8���{$���\3�8H�2I�EÙ;dT�с@�ʓ�!�**��m��Xw)�nh�a�e_9eM���^���w�k�;�J�  R?!�Ԩ��v�;D������ j��A(�F�KU���	��Pp֭rv�Z_9A7b���������
�G���:\5� 0DO�-8��%�ت�H�L�
C�����#��[&N�Y�Zjs
ΐ0A>�	Ń$�m �^2>tW��"p������36�TiJ	[�"gP�M,�*yl�{r<�4M����	]+�C>�y=T8ҍ!'���[�'�TDg6�E�
�I��r;q�y"d���iI���[
2,����X��V�.x�'�����\d�a{.z�D'�C��d���7= �I%6R�Dk�����Ai��i#=�34�f��x�>HIbxč�m��7����ԷV�<⦼���A@�c)��@�Q�r�ۈq�m�ykx2��D�O��6�Q}�����'2R�P���V�8C���l�:��t;��6�u�tƋ@���I���&�����Ms����A��VU ���f��8�r�-��7���)ݑ�޲�r #j��խ�Q7���Ӗ�ꔷ$K�Kوƾ��a=�� ��� ,�F�3�E��>Í�!�E�����WN��,p(°1
z��~ S^��cb������3n�t�8��Q�*�fcg����L�HH[%��^x�>���)�mi
�8��BQC\��U�j�=��Tg��L�6��"�6�63J��O�*��:�ͥE�}��K�K�`P���ԵqDJ�P��� oա%�n%v����	1�D�[lEf*+�K���L͓zkm�Q�6������W�M�w�J(q'�D+Ax�m�����<K�89;S���O'g�D�V5�P��"���	�
��̋��>�gޝ��-z�kY�[��6�Y��-5g� �D��
2����Xgr�'�)�R�W����n�����o�4Z�J�|�n}�ngyA/坯�!>
;�j�m�׃̀X��Ĥ(>@�����ٶd6?�8�J��M$P,�b�_PL6R��FW���-��AV����n��٘J�;�����_��e��.%����*�V�;d�X��P�r���d�V���c'���ML��Vvp!l�e��&��ۙ 'Mο\z��e2ߡ>fҘ�t|��<b��J��)��C1�3^���YF��
��'A��8i�9��J�3š�Gi֍��.��iԿ¸���k\N���)e%��3/Pڀ�P�8Ⱦ��LԱ�
H�z5���t ��0��ԁ�����	���ـֱm�m��l�i*wC�m~�SѠ�Ka�I���14�`�׀L��f��"�|�?������%*�K ����F�o�0D�_��DtF�1��_ۄ�Pߎ�QS��Yq|oU��Fl�É�Rє��/FP����a@�V���
�֔�p[���Q����if�|�s3��79���ۼ�y�dL~�TU�4�+��6ͻQ���;��!W�"W��/em�kwC%�Q^���+�7ʫ��@�l�����8���?��ܰ&kkexW����zc9L;'�ʆ�E��I�ľ�^�O��_>?pv��ܓ&^�Z�B(�~�L�qx�LA/M�D*yʕ��_�F�٢�#2��O�8L^���8^8��z��~�n
]��d���(�
T��
)R��ӽ��a�b���Y�˫\k���3Ff������^#b��YZ���%	��:O�m�|"�K��?y�	2$�{��#Ir���ʺW�L����e�Z�K�\$H٦@x!�'��{���!�Q�?Z� ��X��jw�����n�Y��='2*����������ȸ����9'.i�#g���U�zQR)�_�L�Jn��Xg��!g�Rw� K{R�"��=#��Ԧ�ᾷ��`%�h��')�#��ʊ KX�xW�lE|���Zd�~��S��e�M�Yn�o�#��Hu�e dMfe-�T���{[걜���~s�в��4�\�%m�rod�[3qߴS��g��-��p�[qZ}١m�3b\�+
�&��h"���	����]Z��S��b=����]��,����>#��%��L���*������͂l����V�c�J�r��{[&҂@uܜ�&��+��S&�!7&��b���բ@�Y3��1�����p�ҿ��
o�A%�lS�e�W�ؘ�{ q�8L.�^� �L�%�x-@�x��Yə!�L�vڛO5+�B����6d�b��<��x��7�k���ؒ}�h7�r5/�0���HW�+G�ۭ��ْ��`�LR�!F�2�
'�2���Q`-^�x
W�B=��s�C�"�����I�������8"�jQ��t�(����MyJM�\]�Ƽ���o:�d�0�����1j��b6�<гe��LlR���.H�����I�2�(��cx�o�@��l8�4t�N�l��Tpt9�Q!����A�|�H�&TY�iV��ܢJ;x�����s��Ҙ�e�sr�>*Id��f�_���2�Ih���ީ��G*�?�ۿ�;θ��yj\�D��J"xټ��T�^����Eb�U<6��*I�(A��(�9�?�!�����^X��@p��:I� �j�.�cK�4f�����k��^��?+�@<AS��W`E��LJ���*,�]�dkv;h�Q��S�.W�˪��ۇ��G���M�|�gq:>���	'�����}T�Rg���w���t�u���~������n���^�ےT�h��Xk��o�Ɠ�� ��j6x��LP�q,9Ly� ���t>�uH*���C������k�׊�zB�`�c������R�q��U���&��h�ǭ��,�����������~�K�j��l!�~Ur�#:��sZ.��fn�������Ѽ��L��<Ȯ��ٟ�*�-`�����_s���Ǽ������{�@��L�4�VZ�ƻw��ϐa% �u����� d�V��͋rY�|Q#���T���8C&ޔ\�Iӆhᚅ��!���S��:�+��˰��L�c��SiG
��S���%�f��y��Ґ��^���zB��$���ɼjO���C�+#�$��J���7ǽ���X�4�6y]��~�˿��N[99d���[������md��$��@��PѼ�z�?��,ŕE�^��E�-�<e27�@r:�1$Ejp�NE[f�T�l1��2P����V����P�h<�$�H6�iM���V$ӯ_���*���X��,�Y$�3^�l����^4j�v�|�g�2mT��E��ѠߠL�Lo\�0*P����o�{ �\O�q���6�M8�Eo܏9����>�����aQw9��� j�h3�{����� �ZR�o��6v~��:e�q^M��@���m^@d��$|��A��֜�̗���m���%/�VM0��u���PԱa��ͬ/��Md/�.� 5�z�n�a'9b�#,GY�W ��ٰ,�hF�ӯ���iD����^���A�}�bv�lX�D�u��/L�I~ >
���q��SU>����Se`�C�H�r��
��OYc:+Zٲ�n=9==��n��<�������*�Ւi%�zL�����fk��B^�8u��t��~��H���LQNvSX�PQ�S����fa��@��ˏ�dÏz�C�ŹPd�ɗ  �~
��Mr��h���d֘���6�N�9:��,+�SM���<�ƶ6����&���d�Jϋ��B5G�\:ӎ�������ac�Ҿ��U����r��$sF�� ��d�̑V0c�F ��X��y�b:���$T4I )"J���/F�ã�L�U�6(��"��e�N�\����($
EHC���Wl��P��3�!2!@]�l :��A�BY�L�OY,
��F-ޑ�Aa�#I@)�s��r���!7�C� ve� ���!�����U��rEÑ�AՆ�9�@u0-JԅXB�J����U(�^ �fV+��<[Λ�)v~�W`��g��,S��@�PeT�  ()IDAT��C�@�"���<�k����r8:����..;��x�p���)=�p����C���$�ͬ��e9�%�t��ł��*o�[�֜�44B.8u��o_¯W0VsW�7�]��0XaƋ��N�
�o���z������(�P�E����@,��K��dN'��^cn�`H�X��L����F��<"�Y�]�k��
�eb(Җb�TD֠1�=�-yc� �ۏ@+~[bc|�3n���@�y*���VgQRV�[��[�E���LS��Xu��1�7퇞�8���2�	�*�B8�Ӡ0��i�����;������	"���4�bh`ű�ULy��]>���}
������)3J� �`ZuV�aCwO3g�)�~`�A�2�'�
Oe��-�]����M�nG\0
�=0P��op�s����R���k��es�
���j�&���<H"�"	%���%�W�S�d�y�d�c��e��6��i1o�\e+���T����p:��l�O�=�+ZK�*��t�s��J�^��H��&�)��q�M!����#�6����H7z�BZOm#�e���̯�&8���Hh3u#$��@Qjȥ?�,e��P'�?qѴ��ˎ,����C��c����s:$���&w�$|˄J�h����ɣ�1�fV2Mg易�m�+V��K�1ô3R�b���Is~U~����p�������<�1��јr7���)��Y��r�� x�Ϊ�8/5�r)�FE(\�p6�� %���MHje1
��\5"/l	��5Dz�9�l��Df�KC��x?�� �� ����N��B%�x�"+m(�'�x7xU˪W���R�͂lK���$�خ��rk��3���0״�S�L��p��~��f!��\�PBl�V�f2�WDE��@$E�wv%H"yx6w[$i��5���@ ������@��6s#�x6�mD��[��2�)�9��iW�T# lI ��2:.Ǉ0U� ��3��3��S��%�1쓂�p�˛����Hɷ�a��9�{h+�����r����D�8�`���:1�F��H����������uU]�e0�64�j�Q<�Jqm�-�0���q�)k�k�#���dj=F��X�#B�W��q�˿)�].iW]�GXM��F��*,�<e����б��b]Lx�WF|6�3���&IW$�P�Jɦ3��;�<gj����Q7Ë.��E�5�YFD@��	�eH�2/�8urBB�?Z�b���#�ž���2�.sx\�-]�V3qKoUc�1~�E0��(��C�"FF x>��+1M҉����^c]�Z{��^��͘�}�2[�8��427+�ӡ�$��j1G$N	GuQ��jH����7�cDdB8(�Oe/�j-LP+�]��b����4�1��<T9��~Z��<�`�R� ��;�^G�?�Ә�$ֵ�.(���,�U���B����u�ԚX1/&vM�`��Ŭ9X<۝Ъ� �W��0hQdݭ��nQ>f��߳��h�����.2��j���M"�������ӭ~��������Rd���ˇTQ{�m�3�ҍ��O�mT��=7�k���Y��.Qx4��;�W2���o�>����c�-N!����%��%�5��4+p�YVىB�b�����% ��ߞ	Y4D������Z�$c��g:�R�^US���ꮤ�/ioX����=c��%!�b4�h��>ς��5J�����X�@���=��A�f���d]f�!��8V�%�w8��`�R��_;�*x�bWī]j�����v��ǹ�;�aN�5�:73�x�U�2������n?
B�� D0a�[ ��<��L3II�h݌X D�4%�m��%�E���ީUϊ
$]����u/���/��5�?���	sZ��)�.�47� Di�PY>�a�v�b�-�Bh�r�l�M��Ѩ�Ǌ`B�.�i�x���
�͑���_�h8c�#9a�0�9<�3r|�v��6��ؗ�nѿS*��ڋ��5�|߄�Е�P\uh�NΆ��-�0�JJ�u�ç\$�%�Ɛ���L�d�+/��	D�$`	d�4�&P�T�r�@l�DWۓC�� ���!����s��o�+t�O)�Е��8�n�Y/�(	e=�nG��I�����gv��L���4�F[�Ft�Ӻ�Ҭ���8w�ݕ�[ u�l,&�M�_��䡕M,�܅�5��S1 wٻ@䰪-����Q"��Ȳ�ؐQ$�1$��3�C<�kjT3��]�8h��ڔ�W�Ȋ�,^�R�F��YrT�'s�Tr�k��Hb��a�l���y1|�@O����g���R�㭍���{v�nd*�$�A���k���l_��-������س�q�~��q���2�s� ��p�v��c���?溊V�x�m؋��}�!��SF�z���B;P�rO�����OS��(jS�����Ⰸi���������I�1<{�{�z�r��C�Y�g+SC��*lEH�� 5���=�AGLii�ڑ*�tzZ���T\W4G�׃	K�r�{6��A�Q�U���;����?���?D��睷�!B=U�#�����b�/7�K((s�Jx��18�u2NE�Ĭ7=�֒	6鼮��5�!��wA%Sɔ&�c�9�u�>G>��H}��I�(D�����Ξ�9S�:�zn6y��0Ҝ�Up&��('d�N�7ru6qe ����}���Y,�K��5X��*�h�%�2��w�a��rS��1�sK�f)ڟR
&~	$	 A��*�%Ͳz���D��Lzm�^� �V<�e�B.�[��+��z&����م�PYcAܮ���5-ӟΡe%�g6G%YTW�tz U0��\s���sn�G���O|�B^ȼ<�N��r��b������w��6�a��Q�fez�o�j8C3r��!���4E��%��O��~Y>>�jaBQ��@Q�: ���Ĩ�̠GS"	��� �-+����ԁ�n�1�0Gl�J��d�C�Ч����/�����J���Э1#�F�
+�oC�T*��N�@�*�hheU#�)(�;��^��s���AFb�Ɋ��pj�m$�*�R�Z�R��jG5��0�s���s,�zX�7�^�S� ˢ����ec=54�xƖ���G��Ţ|�d���
��&K	hĉ�d�ɤ��N�o��21��m ���ռ0������:)���M��=:;�oP-A��p)H�i��0+kR�+ow����=$�:�u�֘���윾�楘��!l�P���f�� m���V���u��bs�6�0�T��2EӸZ��S�*��V�,µ]���#��,glw3E�	O�X�&M�d�#/�i?%Rn,𷡥hT8�F��F $x#*!�vD����*��u�n����H�l9��^���Fbt-��V�m=.�e�i-�,���Y3�^&�:@��� ,ͥ���1L�ٔ+N�+� �rׅ%n����N>�����.�=���_[2�D�W?��s�hr׺�����p� 3��2hK�H��AFF�0rI���i��Q%��}D
L�9�j`!Ҙ1
7�Z����0afML���d�����ɜ��"��z92Q� �, !R�I�{���0{|��#��&c��L@q#��v����� )6���ǌ![]6�e|f:> n4�����m��j3����L�5�9%dE��o�"�*EVRۂ.��8k�U#⥼4�a�8�����s�KOO��"~��+�E��@+�ە�,�>sG�L' hЯ�( ����l�1��9�1E���lfN<P�� Ќ S�6G�.��z@����o~��_~y2M/Ʒ�o������,���_��Y���ړs|r�� ���Z\D�ц|1w��3G���,���4%tM-�Q�mj��G2� #��Nel{�5H}�Y�#"[j����В5%;��HF���3u��,dZ�сT�:#�uJ>R6e�-9x�1/���0�$J�Z� C��E#V�K���&,�ɧ��NDL�>N0sjݣ��^g��p�l|5�X����T����~�( �f�}#r�}����5��p4���ΐ��S�l�N����pZ͎��ٲͧ:�ؼ;U�t��Yi���}����}�yb^��*�e�U�XuL@g�A���`�9��W*.Yt����$�*���� Ҁ��K��r��K�Jl�0=��,����yo՞��Lk�$�
^i��4���A�Ę��X��v:{�){�g%��1�6E^�/�%+-��1y�����ȺG�Y�<�%�V��0 >���)%�xD��ٓ>/�B_�s�����D���0�V�S4�Ę33�A��̨��g䒈j�?g��i�� Z�UZ5֔	��FgK�Tb�k�x�3(t�A d8G�F�A#1��%�!B�I�ѫ� >9�d޴4�f[�e�/����������|�E����'��vm0���@�禭d�s8�r8�{��?��'�|2<88}|\4Jު�
��!%���n���𻜺�������Φ�%5���¥h2g��Ja�Θ��DJ���Xh����(������W�C8CGs�'(Sq��	���I�a@���8����w�,B�/�� 2����Ūb7�E��(����LOOϙ¸�i&�h�vK��I���= �}��g_���_��_}��g��j��mg�@x�������ᛯ���O�'����̑���������z�*,@��/�GR�!���΢�X�X�zy����c��6ʦ^�� 	b���Ӕ^��0Q�Ń���H ex1�Č<$ަ2!9:��ƙ��GK��i���-X�^�C�B��vV8�쳯1PUd@pA����ǧ�ə^��q���Z��E�Y�z#��������?cf���W+��#�#J�)sXL޲�:������	`��NoO��BX3ʹQ�[���yw^L�1�����U�y�l&�:-�H�E,`�%����Nt����������Q��6�=�x{�g#na=-�cb��`0�{�.� o/�d�]w&�A��X!ܝ��s���7B6h�x�����ɷ��"�����pQ�9l��2��&�$��mؒ�[��)NGon�S�c9�̢a��@Sӳ8��tz���\u��v�(�293�/Dx�_��5�լ�jWS)�'j"m��K��*�0k�pGt�{��*� 
/��d�����d���p:!)�.gwEH
D�����ߌ0uzqE7bn�FiZ�ѕ�J��ǈ��XN�+�p$��*B-r �V��,=��T`�)P�
jx�K�ʁP~�x�-%�{J�O4�3F�`ʟ�0bB��2VXA�?X�{K���y/�Q���w
xc��q@��@����{�vY��t��4@�,�,	ԛ̥vFl�+�����"�GA���5?��G�z$���As)2��J���J�
w� Çs�i+�W*]r��-�ʩ}X�6|rEBB[$Ղ&��L�e1��,3{1dg$�K$�#�r��E_��!qP��pȘ���V�v��"����Ȟ��7�$f�{'p[�k�3m���R�I�57���S�6��~O3a�v6g U鉉_%��cv����d&9�55'���B�D�Q;R�Y :�C�A�SD���򃙠�L����3`1�g�C��8���@N�X�_��{�[��Y�J�CZ5�����>P9��#�&�gpzhm8�9��%�h�7<�A��[d����?�;\ Q�t7�.��\!R%�	��VsQr$�p1B�&c6nsKL��*[��:�d*�3�t����:U��<&�d�E��m��=��Mo�|�=�Э������F���ƌm��"��n�]��lb�y����o�2�5b��+���EɈ��"��,֊�^4&� s�Eo�ѥ�,�����Fؚ*��ɐ��A�	s�ƭ��2�㹖Y�4a+��yW�s�X,��(#O�x�C�Q��+9+�s�)YPK�<�m�i \sq<�QǏ��a�����W�Aΰ��|����")������l5��I�.Ô�ɚ��'kW��kA�n�i�l�暇+�^.�@��A�5��hO
D$�\$�� #�Q|��sU���]~[�p��Vg��E���+I�Ӳ�p�yv7K�0���!����ב$�V�j+�i�'3\���|0�G�h���3�I	�蔽%��1�qr6�:�y>g�_o�h��p���A�����
�f2�׏Y����vQ���9���8�����.c滮��1����i�v�ӂcl@vtt~ُ�C�qx���+��LC��#{�1�۔!�\<tv�Ϧ�x�0v�v�)�A�!�IPD�0y8�گ:=�q����b�����ҡ���y�hU6��;��c��9X&�8D�I
�-��ŋw��?�o�5xL'�g�R�H�'j�*�GO��O���[w�/2��>�{̳�ٵ���qy:��r ����f�����{�A]�����FWᬎ��7�l9�c�y�Gp�}��[R^
��K�B J�#����互gH5�J�0R���|k������Dd�%�S(ۚǒ�
����p ����2���lvM�) #�Ca%�f�<~m|Ge	�+`�(�}IYjD��LS��B#E<�U���պ�L�"��]��oH�.�'A�#,�0�U���F&���Vj�3��Չ%�򀛍G�8��k<�FW�ф�|������H����@F.̹!!)�g{�>-��qM���.�lD���&s<�Ҕ3��}���cg�l��/�pe�>�e�p����B��?XMwm-I9�������	2͋j�B@r���|U��PB��_\�.�k�&Oze����;�cF�X��GL�O;��q��f���PU���b�qAh�z],h�'�^|��8�԰f�k@��5�{뭷0�b�=�2J����*��kʈ8Kɽ��g� �y%@g)� Kȳ=n�6us�}���zД�M�76�+�c��x�=�z�V���.�3�� 'k������{�C��5_�M�~P�n}(���k��-.����cmc7E�\�����@]j+��L^���Q�&�9���X��-����i�҄j�_�0����WCLu���@F��E�3�`#�!�GejWk^n�e�����b�� 1�=��F3�0���;x���;�������Ғ�vC
G��#����uڭ~WId�����=�Z�vz]`㊲�.Zy�[|P`�$�9P#�	q�R)�<nL���&P��̪#��f���
H-S��x��NИsș%�ʓ�S�YrU|G�V��+�#����=7d����_g8��� �9x�_��Ȱ���v�Nµ�v�<�b&���.����M�Q��9�1I�I��z�O�(�����l�`fz
��W���k�"
h8�������	5/K��G��d
�A�k��ό����IfO��e+�2s�bO�l(T�ց0��@ ������A�MZ����o:!W	��V���xe����F�/�]F��a�.(Y�Ӡ���8L��׀u����9h�x�/���h�E<����s\q�?�%��?���-�\��^dd�>|U�k@�@.��8�E�Wҟ�~���i!]|f��"gD�mpt:�.���,GJ���d�+Jx���a��ɍ��,���KlLy��LeYW�p���\8�$#��iG���7d��@�DZ�M&�Fy}d�U$C^��n��J���Q��-@z���gi�����:�Ⱥ ;H�c�����Գ���Z�<�S�\s�1~d8���j
`1��o�3XD?�yF�� �x�t3I��'�@���@(P�%�R`�~�
j��T�ʨmb��`���}L���[b���Yl�t�Χu'�ٲ 2�?��w�����7�@=^;QI�ٕ���u(J	��j؂f'%�`�*�O`'4�d�Q�t����ń^��2ݭ�r<��L�3I�$q�sE�4:Q~��
i��vC�����(C��p+�5�|���d�xJ%Y���~��c>P��=6jj��Hi�]��8c �w����/����v"g\��P|�?�\��]$!>�Ii/�,��TB/&�>gj����3����>-�"�ukȩelKD��{�n�[������@����u���RHzoG��0�5�A�ऑ
kE4Sb����&T��Om�R/�����Z��F[�b�.�^~La�:H�3|��0=����7`�vy���[��lQ27��5�(����ӯ����ｓ�3z���(lw����O4l����a<دv�q~��p�� �l2�p�[a{1�d��IxOE\��y�� ��y��;� N�G�z�V��X@�⎴�{`1f��5��aW5��M]舒۪e1��Ho��*�f��b��lg��7�����%�n�7Ϟ�p>������}��>�C��S�a�HV�܌<M"T<���&���@63Ѡ8��e\�P�z�zD6���S��.�G����t�>��䀃�3&�Z����'S,06������f�����{�Y���IF3�B�#�f&����:�@��?W(�\��Ç�(G��-��A������d���%����1 X�I��Λ~����'��>�5WTq.��	�XL�3i�1�2�^?��G�bm5��1�Bӻsg�*��iw~�%S�G��޷��_��'�*?z-� �-�Adx�5��T�/6o�A$&6��>Wh檱D���@�zIƅ{�������5�կ���S����OQF��t�V���������x��?��g_e�����Ī�5@��@wS̘�R�%� kƿ_	O�*|�;�"�*l/�۹"�`<�����s= � �m���j�:Yy@�����A.�Bty剿Qy�}��~O;�w�q�t�fh":j��ڊU&^�l��l�1�X�Fj%*�*��g�s�u��y����������>?`��
�H2S�b9�!	3�4�&�6�?r��ԑ�*(��-��m.�R��]�4:�p�����_�F�r>{�6_��e���W�$��T9>�^�'��o��q��U�Q1�D�~��!ky� =k�������m�I�u��%����r%�<��� ˝׈Q$�������닃̉�R�ׇ�x������O}�'=��w&��d��h�t%T�M}15��V3^����ۿ{x4�{��(N�%�Pg�������Ϫ������������O��5��.Ѓ�rn�F��P�_���3�d�3Ig�/�:�lHMo���1����ޛ�������{�|�������2v2��^�`t���ν7:�Yst��s��7;�Nm�tT��h����MhP�Z	5�(;�tbZ#�k"o��w#��/�x�.��t�����{	��&����`U�Z�1�1�,ڼ+��]�����7_���d�rQ�4�bv�ٜq�E���������������o�(�y"���%saDfRǰ�Ҭ�z��5�/yF'�X; [{[���˲3)�<(��@�[��}ʗ��b�4z���_�u?�X���w΃Gc�U�}Y���[E ��D��*��$�Ցb�s�![=/	d��$O8(��\�F��	��L�m�n�`a��?h`4�d�a��$Hd�U#&1��E%Dd�ਗa�p��EC^�L�^��ՠ^Y�*6aQ��ٲ.�Yx�^\��ΰǼ,��7�9�2���|�a7����?�@R��:��
Qܻ[�!��4;����1����Oc>/�.c��q�+�f3?1B-�B ڀ֔��9J���ɛ|��1ԋe�9��IepE�%}{T�1ǜ%KJh>��c)�M-�~1g�7u�	Ӿ�����ʧ��5�FgC�Z����wd�{��ǁTuʡ
�0p"�l�c�Q,N-�i[�|�v�>�f�y-a�BgP��MsQ]�G�s�4|iN�&����1��{�_��0)OKh����* ۜsB^��dA�b�ۀT��ڣ$a����R��#V�����p�� o$8�aE��w�d^C���@v��]����}�����
���Ȯ�A������̚�9��    IEND�B`�PK   ��W��(��� _� /   images/b4c55bd8-374e-45a4-aecf-ab43f4af1abc.pngl�tfA�-�Ŷm'�/�m۶�_l۶mv��͎�t:6:����s�}�W{T�ZkϹ��=��(eE)$x|x  �$#-�
 �a���a���e�w��&07U)Q@�,��?��B[�RA@�φ@�� ��� ��P�e �`��6������?# �_���@��������߿�f�h�ff�l�����_����W���`��;��2��',�����u� �o��`�2!��)umwmy^3'�o&�N��@���~�?���݄�`��� �/�?�?afr�����	�k+(��9�Z�r~~����[�K���'@n�������9���#�����������������nbrt���$�+�����������#�|S'wr����w���m,��J�n�#�@���af�d����S����8�7I�������W�����v��)A~��O������W������U���^��>P~����3�_������S\A���uP��ǅ� �0@F\Dv��������ļ(�8_�^LJ�j'�za*�a���`(�����UML��hM&O�2�x��v�]�]���ˑ��j�>�w���ϕ�u������IM�4F�]�����1�|+f�j�'�:t����2ѝZ�&��G-��,	��N]�=<����]�c������>��jª[����O�р/o�s<�z�w��E��4C��'N^�Q֕E���`3����ڽg[��=��	=_���������Y�7�h2t�T�vm�����.��������,���gNܬ*���gz�y�ǰ�OS�Q��vӻ���т<��
!�_:�80?Mv����꣥େE�B�Z��!`~Cw�p�����PM�m&�(|�&����X=
ġ@iTs뱜7�����6����λ����ѷ>(�^9�����Է��������&������dt�l�o�: =)>&:����^����?Yb�$��Z�h#G����m��<���ϔ3�a%����}پ���ug� E)e�x�*W��/!+=yD���5		E�Do�w�nuy_ 4�R{ڬ�$��X$�'+N��eCW�KY�/�d�`�eJ-0�W�qtE�:�5�O["�SBfů}<^��=��c�#nn�K���}��f�x	��z�U&�sAٹ���7���s�y�Ss�\;�z.Q�8��oy�ըB�h���"eSE�����H5v�G�v�UU��\�¬��m�TХ��S�M���U������������7�o&�h�^�3��.N����N�Z��o�*�g$�o\V�%���;��y��I�Q��F	g�!�BO��Q�y��`�YbU�J�$��*Fp;7ڱ���J���`�.�?���������s7���6c�!��C���]U����p���D�n�����$���4���. ��qY�l#	eơ�r�ڞ�3������a����mvv6 Ty�&���^�q:p�Oܖ����r�/�*�݂4�wx�R}7]�[#^6{,�gn[�نb�l|����Zr*�H��C�N�Gx���R�b��3*�Dm�[]z�2&9�I:<��LH!��~�$R�5�*�����Q��n��p84[�
Ɔ��X6e,�7H3�I��.Ņ����~����g'F<�_�p�}���y���*�1n|�/q̈oC��'}���6�=���D	P�^Pz:6.n����FN��tȕޥ-ǥ��R���e�W2�ܖG4<�W���9�(�Ίf�O�K$��[Ж�ƈ�/ߟ�#������˼4ږ�4��'7�w����k܋ޯ޵�t6/I"v�E���������[��8z���[S*��~�v*ns�T���g��1�2�=Uj���#$�H�����v�|ם�]i"ԩ|n�s�,FY}�c=A���7C�M�	q�3kQ_��x�����X 4���d$14�\��sch�ɧG�:�E��g<�3�GU2���`�P�
5T2IU�S#>��6q��˪�1�6M�lלwx�L{+W�|�🰥�����?�QP�C�- I�Ӳ/���q��^�"�=�ˏ[ר>�?�ZW��-�m��Uiٴ�C{R��|w�TN�Q5n/���4�.c�2�����i��[�yE�����{d�����RtʔT0G��G�0�]!�Hwa����8�U���H�F��r�GF����?���&d���+J ]
����6��hic@	���0�2Tgg*ǆU�L�iY�̠�6�V�Z�Gj�q������	�~��י��ń��UK�%�I��?�YY󝴌��\�%�_Iά�p~>K�xܰ�*3.�g��C�	4�����c�����èM&����Gt���uT�ԣ��֐[
^x�1i)4�,��hҦ]��zoç��ջ�?7���[�⻖�1d��x�ǝ�/N*��Vhw* ?����oC}�l��&������p,\S�L�*[��_��BZ��5}.�[�Y�n�~_	z%��w�����D�0�4�4�+�]���\+��!b�sy<b	ȯ��Flj¹��>�>�a�X�.tx��='y�^s�Q	���݋A"%�%������:�?��"�l]7Y�Ȍ��_<�I���C�#�*%��D�Ȩ��Y\5L���nSHZS����CүF�_���5�ځ�F���ܢ�ud��j�0�Cl�J:D�2A�7���"������y�v�A�Y�U�D��z$��]eS<c��Z�<�
��*�"�h���m���tD/x9���]�����v�����O��'8ݥ�3{���iV쇆lj������j������h���"�T3����1 ���y+������{���׬4�x�l��>��k��X36$��t�g�I��X�AYV���ߘ%w'�	GՉݖ�T�����ĉ"@�E������Gj4��M��>��nP�+~+���9{�����nȝ�4�,��Q^pESMIkc8���k�j:�|E��܃�Fu�e�f5�����%��hqċ�;�6��uR��Qp�A�E\NM8b�6��BoRh����wpWxВ���`�o�XR�b���O�&bF�� y��F���1�v��$�<�&�wRyn.$�@���W��������BS4�ꉿ/iĵ��A�gv��4
MG|ƌf�J�H{�N��R��])7�R3��Qס�T3��,z�wFT�d�0/����^_B���`��}p:�]�v���f�総 �Eݑ�r9E��m
d7�o��/xދ�<�IhS�����٘�G����.��6F8@i������N^7y�
.�R�%�^!�Q9�G�b�>V�ʊcG��"<���1�����c����|�d��*S�-5�Z��ڏ����N���,���{`|�#�8?���Q��蝷Y�^xW�WL7~_ޏ��(�	�2�apw :����XgA�w��3��"M/Ŵk��oJ
n��Q�p�V^�X�75v+��/d��a�/}��kS@%a�I���q��:c���a)��H~`l���C t��1/��Z���ffseC��,�J�}O�����L"�1X�ty���k�hL���ʭ�`\��-��P�m��lf	 �72QjH{+�,{4G�L��j�j�8Y�?�;��=��,n��+>�#WNO�?�F	���?�C��.�j������n�F���[_H5�J%�\�E7+��[����"?������~���{;V�D�:5q�ƭ�F�N��No)u�b�Q�-h��=�P�䛭�"~xm���8��fƟ(9�e�Th���}���D�2��!�Dȗ�=���=D��Z��b��k��Uf�l*����gg����1|Sj��!�������&
?���SL�>+��f7�$�����aY��/Z�&�@����	��=?����Z�������d��3��O3{�̃�O0�3%Y5M�z˻�Dj;�U񽗫Z���
��Ac��ٶ��4��k���	���\b�3-��}�V6��/�%���,�c0m-��ր*�V���G�̾簹YY~s���k�>�_�����=�=3*&Ô֏mtc��y�Q�IC&B?�x�G��l*�ym�jӞ<o��G��x\�6��<^S�زk2ݨ���Gk���f�T2Q9Ac�ȇ��~H0�;���=P0]H<L�\F�Ǘ}QA��w	A��w�3սR'�x���7�SA;I0�ȩsͪ�6�-�J�.��
��wE�k������
�2]}��̵��8�C�q?!���fS�����^�=|#��%���mF��<S+%$m	,t�����h܃�!_���Mc��цL���[��X���f�q���
#Fh�f�وȠ�$��y5ܾB"�����,�*�أ��TIT��fn�/
��?�����J��ߺXin�_}.?aH�Ův�z�ue$���_�n���S�b6��@B��HI�᝘�D�����تRL���&�)����\�̇ͦ`���~׳m�˂M��p��w�	�d��F�E�'UNN˴\R�p �4���aa��L��z1�0��N��yom���
$���x�k��J������E��9m�Ʃe3lT�D%�M���5��Ĉ�:�4�,�˳"$޶�K��o����o�Y�{����UD�s��8=�e��B�Mg).:%�O���"����wJ^׺��m�60/���y&�E��{ڶ���y�)�U�O�;,xD�<�W�ϔ�7�`^a�j4��1B�ʼ��cFM/���%h͞�Z�Z�x=�VQ������2��M���,]��j�01��\P*���VX��7n=5�d\++�h��e�h:��]��;q�Iq� ��7_v��>=w1|���_U�)B�7dg4I��$���v��>
Na�]�VdI$/*;�Lw?_i��ۤ��Kû���&Z�S%�7�*�,j~�*{r�Z?3��b�:�q��`o�1N�ܣW�fX��:�	�̕���@�;( i��aUP���z7�8$#��� ��f�u�T�;L?�1 S �$~	�}HoX���<0Ga%53\ˠ]�m�RއO�	�<N���8�x�>h\A�z}��	I��D-}&q95C544���n*�u�rX,�E͚���o��r���a}��ߝ���)�e�QeV��s�Fz'9.[d_堙5�V	���r����CJ���d"vg��#w]����D�q�P��\��⽵ñ2*�L1��6y��E���i����Y��c���H���������B���a؞�����0�=��3�b�S,����zyq=���C�ZK�.2�5W��{��}��~�TI%�C���諾(��O_�m��?íX�\�.
C�~'�cDp����E���_��"�h��M�����Z���Ѱp;�K#RRj=�圚	�A�h�O���1@&DB��$���*}������d�C{�Cr��w3N�&��h+	>c�_��9�N�嗌�A��sIf�x�;Ƹ��`J�/��������93�)B���47!�k�� �+=s���*��\Tvm'MN0�BX��ֿ�zk�F�Wk�Xs�{�J`	�&�2.+iQ��CA�'RH	mn���xh6�~��^/�0�j]X2�vD�pΣl����mL�v�����D8 �.b��m��(hv	�>�t8&�ܴz-O�6j-�H�񲮢"@�f����A��E�����ѫsy�{y�����{�9D�/'�wF����"�D��n���d)\�O��A^�
�x(NX﯆a��֟�`�Ncw��A��(���L}��a`9��G�Zo&t���e�FH�qwzY��I�{����¼+�w�DG�ا7<��lݚ>}7(�����ӱ �o��
�Oxt�w_LJj���$_	�O�i���6	MЩ)��އ��u׫����el������Q���PZ���_}��=۶���4O�=k���[i@���2~i2�;��Ȱ;T�Ue��=`E\����Hg��#�u���O��Q�����7�6q�B�<Ԏ�;�n�,T)3�����N�����6Q�o1�|LR��M>�����P�Nt�9�U�A���Y�������z*֍�y	���>��������@ #ԕ��s�u,��,$�F�|��I����Ï�-������@�$/�Ly���8����L��5Y�L�kʷ��>溓��X�$F�sA�U� ZLbTǾ|�CULR#�s��+��� -�&�C;a�C����ɸ�@amS/Xꄠ����T�]�J���[����44 N��U���koca�����q ��_+HPT���']R���h$�T<�nOW��s�3�);�^���!�s�ՠ��ŹH��G&z��s���Y�������c�\��ZDP���-�Y�����9'\9c����`C�vȁ�����'/��5�)��(�Eʼ������5�6nP��8R�o�
���ky�[�u�Gv	8�(|�L�B<ʴ�� t�v�(���ưϴ@��C���>'�ڰ�9�!0�;�L��J9|�<˶� xaƆ��R��%/x�m����8�x��ZS��蘙��Q�
�<�@F���1��#ɖ ��3W0)�Q����"�.<�ޥ[������C��V���3{�7:����>��S�n d�U�L�M���o���U(,�֠�4��@��:��b&��V�w�-��v��2u):���,T6��	f\;���y*$ 7���� 4bЎY�PR�
�B�
>�{���]��N��C�+1~����0����9��cú#7���*g�f ^YI��!��<�;�DS�yfǂIq�
��fb,_�����O�+���n��tY�i}d�5<��&��>7t,�)���߷l���T�j&~s�uʩetގtv.D�]Ѿ��П����~��pX�e���o�k�1�`���({�C�<h�y3D`�/�67k���e�����>��|e�Ԋ7�]����W�5��.��|�!5�اN`���b1��{ܳ`�\���4F�
�,GG�4���-߲�8��l��E���,��S�S��P�J1�]��n�N�un�_��}���j�C�A�r���Iq�	I�K�ʂxJ��/Y|���{��͗��'�b�d�ԃ���y6��W�n��n���?X}=�,~���������G"ʶ��i$��y�p�$�F���D.�����S�bpcx1�t.B���t�᪑/�wo�{�^�G#���R���px�Qt|�<f�4R%�O�����.h���&L)^�x��Ȋ���(QcU���H�� bKAJ��R����b�,}��-i`�v��H:*A��`���;�p���0�ˣ�V��{5{p\{�B�][w�6��]������.�2�@"K���u>×H���3�ؕ���HZm
-Z�l:�˚��?���9�U�ڎ ��ҳ%��Ԕ�A�#���\ql���)	�¯tS{i��>����ߩz�����t�4�NWr2����O�4y(�V3~ <�4D0C)i�,w�j���7'��&5��oP�l�g�K�j�9L��6���sc�f�ЂW��S�]���p���th昑��Д�h�!�.�����	�h�R[f�;���!�&�zL�L��B�	��uc�M&�K	���'��h޽w&?�2�٘�W����#1�?��'8oZ���:�4P�Q꛾����?ʶ��tn�������PPt@����=e)-��|�M�+U;�	����ڙ���Bxd�6�?`O36u�ť2��������?�ES<�P-�oPŕ����BYC}���� KA�� ����;)ͬ>�`|�>�<�~��E�7So�<�y�i�j��X^�]�\��]�����g�)&�2�q�{����`KњIZk|�����6��k����૤Xy͝dU�&Q�-�C_� ;�0d�n�&�B�*��+�OK5�mba�Fd,��k=�J�D�iBM��SL�ܘ�+.ޓ�x�j>�Ɩ�7F3L	��o�o
���W\um#�=2n��5rV�@<�=_�4������(�Ԡ�c� ���vw��u�p��ጳR�dM�]����J��pF\Z_�<)�~t{���x���mј�f�wAQ�I��AȀ��g+��9tO	/�J���2��c�km0gh���������nޡ�6������	��NϼmI1��w�֤^8&ٍ���s����UBI`[����w3c||��:��#��K��9E�6�\� �$��h����^-P'�GU��`n�1iY����{��
�ϼc�>=�#I#:���@z�
�k�����X����F���y��m���5H�T�IUnɿsf�M0�����I�w^;Vw^E��L�kx��[ۼRe���g����`J���xq��6��ۆ�],�E�fC�� ~My��K<��k%����p,f���	aB5=}�w��v����E��A�V�S������#0N�4p\��璝h�Ӧx�Y��P/���8��Y�Kv��G�����=�����P��.����GH����3I��x�Nz�>�ev���Kҟ�c���=�
�w�e��L'ѭ�����@??�q��oϟO��f�U]߷!tݮb��[���V/�휆1TvFX�4���l�Y����~Opf�V��2�]���j��Wx@�l
��R�tR*�|���k=?+�+6��=�1���>���\Bm�{Q�T���o^�g|ȌyR�BT-|�'�j��5�Cm21q�d�Z`zT+%}q�_�J�(p-�h@���mY߭r}�.Ī
��5N���÷}��g�*l.�����~��&�E�z��z�+Vq��`3� >�z��=Hpd \Ð��b����N7�s�8��3�Ǖ��q[VD��X����QHEy��2Yϕ�
�����1���C�����e�L��
��{�NNG:Z�f+�f��jp,�}n�#/ݦYnbgl�Gd�m`���Ñ�����l!�ot�E��-���|Y2Y����r�{~0Pl<���I�Bl��&�0���s�Zd�v���" ��O���@����T��l�-�b���dqaS��9s2�a���`7a�/��7P�f��4)͎6����"��+�����]kDt4���~��m�[E�xpR�S��K�3/�b�7��?���9���oC	h㔛�����X�{�Lbƈ���q��TA��N��*hK�ɸ<�D�����C�_�s]JB�ؾv��I��P�N#���eL��k���h�VT��|�?�g[L�c��z�_�眛\�����!�~��I���-h�x{2\��m��@bq<'����*�>��>��`���>�	?�Ó%�0�*����DM��:��i!rP�+��Q1k�MY��_��f륝��
�B�
k��T��rk�ћ;riȐV �t5D��Z����;�J�m 4H����e����	Ej�P�\�S=D�hmJ̊�_����*�~4{_k�P4�?z��+I_~�vƨ�}��'6 �B�����ɈΒ���'S""���7�
�}o_����M�ߗ�U1�}:t?c�~�2%c#&o�8��ao_՚�N=�ϣ�9���}���**2����־üo.1\q��-H�ބ�[\+B�\O��&���.p�Ԏjk�I1���X�mQ4�^�+CO<���̖�h;? �
}U�w̐�����j���w��j�c�|�t�q�ç�E�Fs���F�c�=�fӉT��d��5E���8Ð�@�b@��S�sm�Q}�{�]IVFczF�^'}�0����D���T�>����6�+��_2a���7��,�Ҧ��Pu��S�ʝJA2��U�WL,I�*�2]h'b�t ��Y����>a���k��>pYz�a3�y��9�0/O̼Ƕc����X��̧r	VX��S�,�\$�Ve:=q3f?lO �P��+��x.��{؀P*9r2���R>LW�|�m?n��)���o���=&�|s�,�X���=CU|��
�N[����%��CR)(r� ��O������Hۑ>�0LX����~x�D�/ee�!��ޠ���Xc��^r���y��XO��sT�(�b�{n�a�YUwv�L}�l��I�?����TfԞO�P^^�p�Lڢ\FM���ž���ŗzV��aړS�6"�|����U��T�n�-d�X�3^?1��Ñ�2mC_��U��O����
���b2�#�c�����~㣨��nԲ���a?7*�|Nr���;2Z��!�pu=C�|O""gv�2>Wg`� ���XX��G�iLm�Q鸱�T1R,�BY?JI+oC���0	���K��>B�������fG��y��%�r�K��څ]
��\o�B�%�a�4��P3k�#$`�o@�9e�2�,���TV����K�J����,�_�Y�����������E>Bd!R夡RE����u,ߡTt�%�xQi/���X8Љ[|l�ra����1Ͷ��~EU��@�`��AP7qV3��]<ʛ�Z�]�� \�0�VmHF��sJ�+,�\��א�P�>�8u�c/��6̰�P�:V/'�<Ư�k����\� ���$�*�H����:+�^B���%����]>�vG�E��x����n����]�I�3�I��X-�f���:�P1m���U��T����e�!�Fj�}#g.�~�17�H�jC�I�8ȉ�Y����W�k�i�P�	_��K	X�Sŵ ��}� �{�4�.u-�q��� E2����;�G٨���|K��-F��
4"!3�(�n�0v$A��s�:�B�l�[��e�V�ު�/굟�Ȗ�WX����Hm!� ���f�T��3R��àb�h�c��kKdf����'�EkdU��C�Fݧ�'MU�!	�p�0�t،<_-�O��n��R�_��$���Oa33�-�ZX�z6C�s&)��S/�5P��dc�{b�@I�&6*Ǔרb��1j�i��A�9��4����c:�!	,r�H����z���k��V�DP~����5wpV/��B��?�U}ĺ���+\���&EߠI� �(p��2�$%��=GJw@j�2����Ͻ�,����?_��Q��d��[+cQ�E-,� j(���jm8����I��B�/<52(kx�2П2x�3�P5�l����C�:�b�%x�z�����l��A�d��t�vZk�i�c�J��Z����<��&���#�z�BZp��S2m.� �.�f<8�(��6�մ'?o$J��/2��e������Y��8C�d��gx%s)����f ����C� =�f��$�QQͽK���͔�aC��T��	j��g�rT�+[��!;$���x��=i�5�({[��݊�3�\~s;! /iO驃�^�D��A��Лʝ��	�(#+	b�;R���F
LӞٴ��,��.^�CMt�i~�r�������C6�nZy�p+��-d�F���A��4��IV�I�Cy8)_����@[��,�a�j H�̠�-m͛VO��E��[U���AX�R4�4&������D>��&f�-Ӧ�o;C�k�H���e�L\�A�J�k�D���l"zdU_v��DOE:��/4��Bh�,2>?Ƹ˃-,��V꫅����Z�h�E�x�V��N�W[��3.���O�r��	�@n+�BD�`�s����_�w��7��X�h}�!a�|�_����� 59�jG�R>��Y�Gp�b�܃u�O}*�����L���%�尗�b�����Eӯ��`�!��M���}�G���/�{~D�F�R�G�4"�RФ�zM����C����|!��J��e�5Xb���7��7�-0�����l�qԭm��i
��F�iD|)�0ɛ��CmE;7��$S$E��k :QY��#4Nk�6u�)a����_Q���r����9��@�~��v�#��^�W%-�N�̋hUE@�P��3Z7m:�(�┊�Z�
�-�y�~!rO�[聿>�y��>wxJ��d��<���9���G���9��m��l��Q�	K�W}o�߯y=��U��q�+����vlf��b�XTi�&Sר�t%K�_������WV�f��?�W�=�3�	��f�+]Ѷ������w*�@ E��!�/�a�m�T�nE�#_��Ab��z	�Ybm|�[Lj��h���ET�I�D<=�A^���"B@C�>S���X���գ����jfa������k�D��xN6���`f5�%��^B@h$�ru��`���5I����%e��{�2`oC����@ڸ��*O�GA���!�����A�Fp^�3d�Ó���`�N��l�Rl2�
?tg��3=�5�/!��09��kS/ �J/r"s����=M;]Bz�<f�����Bo�ql=���Ĺ"�v$����?s+M�j���kK�ġM���z����w�ۮ�xB,j�{^�g9�֋0��Z0A��ڽd<����-�#e2Z�ZW�V�Ixض�XR��ռmy�m��	�4 ��kh��L�|k��N&��j�;�~���V���k���H�1]�h�t��`ө嘩Q���FDI�z`�"peTs��G�c�����8�I7��ԏ`�	��ta���T��B7'���K�Co��r���=�ݧF�/y�|q��ew@�#�Rb�\��T��_���Gc^k�:><��R�b�{��tW�'��V�(1�&�8����(#�kW)��#cv,ٕ/�����,���5zQ�92��
F�Z�zx?f�����kA
ۦW�4�w����k�s�/�:�J���n�/jûd(iĊ~�?T�kg��_0[`0�8���tQ��R)b�ܢ^ ��M"�}u�ݎ�}��D7���ҫ~��:���rEU�zGZCD=ba*� thP���*�L��J�i�{�yƆ1�$�>J�W R�������W�p�W.J����
_fv��P��j|mq��_��eQqs۩�4E�*�i�%d)�T��y�g&����Y�ZZ���|)�V�Gl 2��3����h>:U�Eod�8=�*n��$p�T�୰��#A���TCbods��t�WG�g����<�*����:l�F/B��������1A�6lR�L��4_,���1í�m��������zˋ~r���ָ�v�ܞV�KdrG�؍LD`B�[љ+�i�Q���^�.��:��&��"U����v���f�έ,!�z;��h�1 �h�N'0g�Si�I���_꾎���;�c�k�m�G����� ���M�"g��v��k��D�*��D��$�TE�b����m^�C`Z�����[���®@n��`n�lQ�k�8���߅a�Ԑ�]@�\ó4�	�z�;�{�D�^�_��R�l&~�呛q��n�����q|{�#3-b��F-D��� �����h���2�>?�6�R�se�])k�z
��ym}�������04I�>N���B��gzCࠤ�i�>��Z���=%��4�R���w�{�K���>��|���_r�]lg���(��|�7C������k���ۈ��6�?p6[���'��}*q��᫯9V������M�pr�<�����m���&�	Ä�HSc� ��aH7��]�eTl��*�KO�x��h�=#v����wɣ�4������11�#):G��~�6p\�:����^,"��21��jC�x�ŊP�te��aܿ�i���\i���&W:�ƞ���S�J����E^_��{,q���5��X<"�+��4m���Н�Y�mޖ�JU�/�ss��O��>@��_���K����(|B�[ta�d"�������?�[qa:�o�hd�bf�~�,�ⱪ�2�Ջ�^�2,���?��0i���g�P#� �����50��v�D턫C��ҖSY��-�y���W�3���I����G6g�!�X#���
�Ʈ�L��!�H�S�}t���tͻI��\*/P9�X�J{���G�TЮ�94E����=�P�8�3D��3����8b���}�9�V���Τ�^�����o��TٛD����;��`ߟk�kb$�b��׷ᐵ���Q�}�_%5��\x#�����r��N�p��� �3�ځ�<+�F	$	��
�op��#�S��{��'�u��;~w0�}|��a�n�FS�ֽœ��s�C"�S�T��r���"Uҵ���szz����t��፭�?���>�L�0H�ɨ���Ă�hũ�x�
)�ħ��)�� @�b}\>u�X�:�HP<�U��V�,���(�MƏ��R�Tr����J$`R~��U]ϙ�ԛ�����nd�9<�2�����ß,��CnK��-�S����n`�/=��6Lď�'�Y(���A��:u���e�+���T�T&�ͧ�ζ�WE�+�j��{��:�P-�LL2�I�m���R;�Ʒ$�B�f��;F��E�ao�b�&Ubol�ǰEAk�wx;d����X͹[���:D�#t�ц���0F��O�YoÞ��Z<U4��={�pb��, �Z�F%�n�ԔO�ۑIw��us[,�J��q�T޺`a��1(�*%�]�K��o��&��v�TDL*k�Y^ݭ���4�8��pl�u�H.�������C}��~���!�jQVK %�Z��$�"8HyU�m����4�-��4�m�r9Y����j����w��*�<�sC ��ѐ�$�z�k��PC�&�M%�o(E�ma��@���}��4�TeM;���r����Db��m�M^U~\I%�}��� �=��Q9~��v0��Dv�K���Ǫd��ego�r�E�JB�"��2/��޶-
�q��i��V��F�J�����d*3H�"`"m��y�W��U��o쫉Ib����ڿm0�9c&m�����_H.�[X�L�2h����1u�n���Tc`�,�gI��T*f�KUРH���f�Ͽ�=����)��~���eiw�&�~Q��i��)��!;>����Hxz���� 
��,e-�Ծ��V|�R�r�1�(<��g��B�O B}<.=n��|8�LB�AZ&h��o����%H�nz��_z���i�|�2��T�<��Y�.L��zSHf~olq+�I�CV��ۊ{��x��j���%�3Ly=!?�h"���W�`�ט��׾*�E�tꇊ�.iYT;7�(D��'M� ���
Fd��T�vs���o�����6�5o<󘤶�4��_U��GE����wި�V�'���9}6#����8����7U���|� ~@�)$��H�ˊ��:�X:P�����Rk��W���;�����z���c�!K{�6�m��x&���N$S��/��Ri�[Nˎկ ���}�k�D��YI��D2�+����=���&�0�rS�]h�X�ԓ�r7����?�R��Z�9D��	�Lx�=�R��v;��庙�����YּX�h���=,�9Q!���"xz���� ��ز�*=FF���l�v���	o�B��(��m��<קT�4<�2ͥ�?hF���iH���ч ���?q��Ә��)�ߦ�1D�qb	s�"� ���O`O�4ʁMZ��y����Y����ȿ)��a61�j��,Q�l8m%��9_��XfnYoy
�=��y��¼�Bo��!��Vh������j��I��&�a���	�`i��2r�a_��m@�+8��fGݿ~Û�eů0�y׾#���7��`ΐ{E3�i�^n�����һ 7�4��țMo�U^�[�����J2�6�46ux���	���BB�,��9U?�H��O��^�/c�~��Q���V1|���Wor��`$a�D�-��o�?n�q��N���9�Y�Z3�1i���.��6��p�R�%4�s�����,L4 ����h=F�+�����.�:l"n�h���1�4K
o"z__�|�����fB2�Ī�[`���>�:'���;��a�S����5��G�Lu�	�;��fgE�ցQ��B{*��v�����s����z)�.k��P;%X]��v�[흜���?��Vsj�rF]���<�xa%��HSe�`z�2�x���b�7`��O�F׆�������yC�-�m���V�pq�UD��\�%x��uq�6����˴��W�6w �ƞ_��F��� �*��ևe��[��i�E�&��M��iщ��l����2V��2���\'��������]�W�g��@�%6T"��v�?����X���s/��s�K1�[1ө
����;g��
��z���G�L)>�T������~cĲ�Y#@V�$�Sb(Ha�eT�����餀��'�c�	�� ��fU��9OGyAw,r N�9y�*Ⅵ_r���:�h;����~�+�7y�x/Uh�)�_(�\CNF�����>q���iB�H�F!��Pb��[B�{R��v�
�S:�W���>���;#��qQ�������M�b�]wu!������j�L����r��\�m�c����mvn��=��`�� �b�A�d�����abM��,�U�����&�9,�ĵ�\D��b�7��tE� �#��ٟY���f�Y	�"�$���/\Q  @ IDAT���#6�O�	��W�:h�u��6k���|�FJqk W����ZvZ����^`ĎLRA�x�^�XM|˵�c':0��2R�dP�^e�Ԧ`��,7O� X2^�������:6	q�d�����~���ˆ��Ri[���$�"�C�~��տ�1K�)l�	�9woY�%�)ʱCsXe��{��x��<��n�:A6
s_	����L��*���:\��6u�h2@>�����m{�G�zX���I�E�:@�(�f�ZBѴ���I�G>�iVM3�,�+3'!p�f�d2�Iڢs����R��Z�ҩ�e�7>w���l���ƣ� �Z,��fm�0K;���m���������oy�X��i�_�=VJ,Rl�̆��v�{��O�O;6�aE�d��k$��Vi��X�v�}�V�#��-�o�a˒1T���촦��9twR��/FX����	x�)�y���o�',^�����2R�`���	;��'���J:gڡǜ�&N�؃������M%"����4�O�� c�﷋�ꊋQ"���Y?��9�;���ɠ��Ѕ͕9VfރD#Z��v�ԋ�8^��I��Sh���آE�(2d�^B��������2h}+��x��?�'e%7X�"��PӞ�:���k�7��g_pݾ��%�X����q��7؃��4��^�14�R&(V��@���Zϣ����I���"h���}��v��`���r�啸� �2��F��w~�*�	̮�^�6N �ؾ���f6P
�
_�k]�-�)֫���駼�����m?��ŭ�ٍ7ވ�]M��p�g�4�Pu��"�Y���
�Fc?��+u�
��P��I�*ƨr=��� |A;�෰I��f�o�����fW��m�/��#��5wZ4I�Z	_� ��k�5�"Q���$m]�'�Te�;Y�7	�X�8�8�e�}'���XE����m��e�K'����-į��o1�� rB��(�8��?��!<KR�U g��.sn�y��;�A���fL��\�b1�5��x�V������ʁ�QaT�F�f�&E���Ƽr����y�+��$�E;�=l;�6�t��t��<�tڳ�P�x�]��_��10<�(8S���<VZ��n-r���'��-8dO���$?�_Ax=B�J%Kz���(���>
ZR጑]��-��~�����$�y��ǘ�(��z��b����Ŕq�q��wۜ�S݆ժ.1�q0��t����S�U���*U�y�|e����`w�>t�.����ż���4���Oħ�=��#(�Z�x޼y�U=�Ү���%�>�z�5{<��S�La#�+��U��SP���D���-ʹ��}�����*?|�#���럽M`L<
X椊� ��V^�KX�'<-*j��ٯkЍ_�O(�&]��XH���[p�w��������rp�Q&n�N.)��i?���ĩI��Y���"@�RՇھ/j�-[��
�Q-RãR(�L���ϣ��Kt���[��=�f�juP��g��1t�'*>���`�L�J��C�1i����~ �w~�������LᇄH�W��U�ɚ�"B���
�k&\ˬ[E�- ɐ�P8e֓dQr!
�<1-�F����$��N��Z�Y�VnL��\��J��9�;H E6C�K6��+����3+6�a��3��(��n�:"���o�I�f�ngx��"�%�U�FA؉�Ximm�['�t���rƧ�b��>�_ml��|�q��#�����I�E_����7Q��~�2�f�!�n�xP _ɐ�V��4/�p&Y�?`�̧��n��A�eM0��Y�=(|pEORy! ��$H��%����: �;���!;��pįv���~�L<^��cAn�>/�����#�,�3�b�Qp��i�"�}���ʝֆ�
(�@L_s�������̻�Yvnw 	��Nn-ڛW��\�^�q�xs��A�Ll1o�aV��)�Y�^�n�.\Su&8�Y?�偎�V��ݏv��V��h=�AQ& �-H�L%�5�-�'�Ү�THՆ��n0�'��wk^�@	r�>�&^����w�pXz��r	�8Z���Q`����q�pKS����bq�#^�R}� �W�YF�.;&Ski�־(�� ںd����5�H� ���S��@	���5Â�\�pS7�G�<�R$�֚4�������~\�:�3�r��-`27t2ϒ�p� <�$����0� 1��4Z�-.�	z-;e���3�ɽ9������
��V�js�l�@� �t�U��s�ҀA«2�c12+nI��6�v����[����ϩ�!���\��З���1x��G@O���O�ڬ<�`4�WF)�@�b?�ǘZ�"B��eps]��R�����#(���1�cvT����	J�I����8� ��&^.m��Qѩ�8��!�̀I��_y-� ���P���V�2Y�I=(l%�p�A���=g!�7�W��khW6���6Q�
X�*�E [�R���s�����]�`����QB1�v�����6��*}hBH��LQ%��EfYO��f�S�,��m�>p��$^�Z`F,+�!@�_�i�2��3��o��43���Z���~p]?�����UĂ)E�E����@�e$Xή��==��C�;q�`�ZO	�����2<�մ�ƭ�����Pİ,�V��%�Y�#���2u0n��K��Ⱥ�����輶!�Ĕ�L�[kl�G!&��io�,)�X���%�NS@<C�jM���#v�_��<���B��rB aN��Hʸ������qw�]DIb}y���G�Ss@���,�~���7��|�z�1���"`9��)�:�|�f��V����Q�Y2hJ��gayc�7)A?]+<2����hr��L�1�}��qυ�2<�wc�8�eAVE?�!A�la�yuxK\_�Y*(o��e���#��,[h������"�׎~�B<�%��'sG%t8V��H�	�1�8��_+��$�'q6�"܆w~��ڇ�N�+
Z��s]��܆0K?5�y��ef�&R��[����E���5�F?�����x%*)e�%��H.Ѥ�4,�Z�6�v��PA`kD��=NE[kB�l��9;*s�I�j� �N��fw~Š�	���B8�`��N��k�W����u1ν^}�Q��/.�s?u�cK1��S��n����*�2�nEY�VC�w	��fSϠ�3JZ�����(�@a��LU �KMկ�}�0����^;zkjQLN#CS�]�I�Q�b\�������X+�C�K��-@1����OHp	�y�l"V�{�bk�dm`�";������jEX/�mk�=���#�*w��1?�C���@�*xS��"E1��<���3�C}�7.T�ҫ2F�� M�n%��p��VQ��)�����곫��2�6���w<�p�'��ax�Z���&FM#)�rO$����T�H����_~��x[Cx�������e:y-���S$��S!�ք)�'�qH�PX��j�N��y�Q&*�"I���S ���'�������>WWC��qZf�KV�Q��2Eq50%y]T1�`>(�l/[L��vh�P���E���~�Ǘx��H��|R�Fzqٲe�)>�{'+���S&��=ژ����0�)�P��l�,�+R|��1�����A'P� 0~��T��L�|���𕢂
��J  Vnڛk(*����#DP�Nn^�4�S/���I	�1��<V�t�K*S�#�HX\G�Uٕh��it�� Q�N�����D!PS�*��O<Ҟ|�	K�M��B)"�`
���0�����)3Gz�}/���I�$( �Є󡚊���R�:��+Mw������5�z�M?b��v51�(�W�uH]Bu��x����-|u���1;�P���q"���Wİ�8k�~��.Ωɜl�y���������1*z8̋/�"A��,�Ug�5�ttLR`uڹ��
�ؽ��	FMm��48
��8^d�����o�}=t�q\�E���8�7] ����}5������N�#z� \�T8��d��C�K��YX�K�n����B����"�3B�2)eV"�u! ��.�خ!=����9jwp3��+*���		KA=����{�ӫЛI�7�+K^�����=7xU�	7Q�l�uE
��圶I��1�r�Zn`��v����T�X�U�a�ՊI��<Z[�M�a?�Q�0�r��nH3Q��7�t�[u��O����9�dW
��d ��$��)-�5"��6�Jk��K���g�p��y00���L����E)1	���W��cg������&7Y,��&N#p�,�3��Q��	��~�F����6W�(5J;QBd��-���y%��*����(������T�����Q��Fyb������o�Ua�	��Kj�yf�Z�6(
U�)�����~g�wjS6nr0�M�攆R�8�<���;%�-��	6��bq��cߒ�)\.��d,"���uQ�v�%���}�=#�~�jX���Y�w�K6L�tLC�j(�A(�����,�#��(��ޘNCxZ#����ޤ��c�Jk����W]n�I�|�ܝP2��E�f��}`n3y���4�g�o�LEm���J\�ص
ũ-���_�����*��܅���昁�Ht��7���#��i�7���a�׿�ͅ��N���퇄lsmk�p
��7{��3�Џ�}��������Q3'�@i>8�*կ�S�>�.���v_�m�^��������daL�Lv��F=y;J��1���s)�4b��8L#ƒ� �e��ʸV��b��J�%�(�(cM��t�V
G����m��c�T�w��J����@�Pt}����<�R�D%)�F?q�!v�z ?�5iW@/|M�s��I[���Y@2�U(���(�����sy��B\�%^�~SmTu�%�m�V��ٻY�9p�C4��煇L��&�y2J��b���[v������Č�ge���9����p�A\�$Dӯ�iXͫcE'XbT�b�m���:��/�z��
�r���Tn��"�@з��n�ߍ���o�A�|Ն�O�c�� �c>�p�%�wc�S�%��n�D�q�(���ږ������v�-�t��^с�x�<9V��_��TV�&,��*�f�G���6�� 5b\#��7S*_�:J��\J�G�7��ģ�`(�`J�0�C̜ �~��΍I@�;Q����ڗn�Y 4�l!v�ʣ�"ӏ��ăA���P/A��w�D���C��-��kS:x��r���E�-o����3ћz�-�O� �֒����B�Bj.���8?��K�b@Ѷ�>`���(�+?�^b�,�������A�%��E�ڽL�T���k"P��N�7rdQj���M��/
L���D���".���<!�  ��]�w��H���]̧Nn�m��M����������g�gc}u��u�g(O	���g)W��֙���V�eS���1�����a���|��9[}�n8v}�^��"���
�-�Q�����~�C�	8
9������X;����Ҩ��q�j�P(5V�W� ��ȏ�a��Ń�ј�m�8�=L�3|�:��!�*����Q\oN�����h턶��"� �%KS�x����At7M�C�IKyh7m��檎�r��X?RU�>W�ת���61�������K4��4�]a	��QA�� U�~����U��9��h�3z��YY���������~wys�=��*� ��&`K�X��]�d�9�%�3�G�!%(K�4�ƺMmO�������ܦg0N����U�S̘���TH���(%dNH�����]WoԶ�]�z�܆g�wƠZ��~�m���fw������E�x���xz�<R�Ԋ�Q'T�'��ͳC`�p1�9�j,��~���*����_��G�i��>���tM�_͆��bX
��ۭ0�O��\j�#���ϳ���)�Q�R5�Ha���ӾN��W"z�&Sބ�ML��٦6�L�&�&���"pX�I/ոhOm+��g�ϙ ն�*B;R���w,t�D�Ƚ�f+=��k<c�:�0�`��:�כOh)P*�%��1��bJ��:K�GI�b�|�	־ev��K*!�"���X�{���ԟ�o���b�)��-�����ӛ����u���h>\)�,w]��J�>̍���ˈ���YkQ����mtV���S?����־׉[;g[�����!��)Jƭ�n��>q\e�$��� ��$�a�e%*�k!�t�i�A*�YO$K+�S�f\ЋO�W4gZ:O���ķEm��R������L����h�t�X���oN���o�4���|�E;t��,�s;�V��	*˭�eݪ��;��b���,"h�aP�\W�K)
�SvG�*��I��`�;n�G{��m�����!"��M��(8ex�>���}�n~�d���<�O��|<!��V�f����jUF��9�uV�{cC���x4~���]�L�j����Y�ɖ�����b����e��y���,)9���@1�O��&k��-$�O���>�M�s\g�xO����,�o(�H�)s;��3��̳��O�?��c���!�_���ݣ��ք����w���v����G����Q��{;e���Ω�ӳ���P�SAK��h�m��a�j\j��UA�ʯ����ۜ.І��L^ +�ot������������,�>�k�n���+�5�%�nJx Jc��_Xt�A�O�	�'���/��V}�Pai��{3X��*@�~ʀ�Ŵ�a���� z�iJ7��Y"��u��W\[�2�].�dq���'U0	������k/���}e�植<~?+��/�b�t�er���S���5(�0�cP����w஼_�8������wdD�7;渓��g�o�W��Ћ"@~+����M���A�Ř�{�}�����k���	p+��玵�gR\$��$N;e��Թ�ߴ���]�0m|s?�=�~l{|�u�m��	�Bm��=W�� N�+s���ÎG�^oN�X���s6�*��7|��{'�����8�\6&�&���I�s�ѱ�������|?��k��L0FG�@��U7×C�+�E��_x���{�pi�@Tճ�� �����L,�\��¬��	摑 <�x�K�w�#��|�Pk�[I���8P!���U�L�H2������S�ߕ�5�N�`y�V�w=a��[#۪T?r/q������.�N[��t(�+7sA!Gx}p��<}�hM���V֎ֵP1b���*��_�c.5K��ZQ~�3J*���=W� ���{����7�m��4~�Th�c�?՜9���u�9!��i��TC��Kgdk���f�!�� �q�R��U��.'�1��
p��}��/��/PV��z���]g}}G������	�l{#4Ìoz�FG\_ǝ# h�)�� Ɲ��G�է���f��I]u\��/�w�r`��P����������"�Opۉ�Sw���ED��i���qC[�E����������nv���oF���xD^y�n��]~uVe�}םY��O�P/Հ�/���'��;kC�U�
���S��9�:��#J8��l8"~T{-Mt�>K�<ְ
y��8�m��g)�ժ�<@�!EI]3?.���
%�����{�[v���鷷�)	�4B'B"�бЋ�A@�D���GQ	<"�
(R�{@��`H�5!�j����~{;����}νw�;�B�H�3�}vY{���]o�9��*͜ OgA֝W�@�L:�+�q.����z���;�'�蕗�j�-а�d��Vs+�&#��!k��4�z���̍��&EV�Aܙ��1~%����)�ф��w�[���$��g��ӣrGl��ii��d��3UB�ɹ�k"Ӓ�(7u����"�}�'��;EM���v6��%Xj�a98GE�,1���r��������}��G�ᚿ�&��gد;��]?����.C-�A�[���f������ݑ!�C0����6��*�Q�i�w���o����� B둼��xӛ�7�r+�����o&�N&9(=���L�cfi�n�C���~6���$�c�l\xZ�t���Lhbպu1���JmT��L8@��"���"���\@�tf�eT�rI�
�\7����K>��S� ��X���W�:��G��8�9X�gW�kR�m1?~��,"F���Ղ�hf�[���FԔ�	��^���/ �br�)�#��$޹͕r���l�<Aq-\�g({�U��{�Cb�{-��C.����p'ߍ2ba���P�M���-g�7�A�5�e��?���$��}��j���>�����9����y:�#x±������k�Hק�p&3���v;VB�y�l�@d�u�N�!I:���t6	Qg���2mt.�Y��.�l89%ε�k�7�vl�dz9�7��q�I��7\��LQ���.���k��\�_��߉�{�?dlcX0�Pn$����=�D�%&2�}�qN�h�N�;8����[�Rё������h6Z�\>f�^���ׁ������%�7@;��D]<�N��,��b��.���-�C\�L ��16r%�&�+Z}T!:"j��РT�kS�F>���/��%u�6=�
�3)ΑD�Y�6���y2���o�n�,^���� �[��]��%�Җ��|��CB+8>���� ���;���c�r�g��!�l��[~;��l�_��;sT%�o�X"W�y�2@c�{:�\�?��Χ��e=�$~�qJ�G�I��5�R���"��Y&5f�dm�K����:�"��继�@D�W�YŢH��Ԡ�m۩��g#����o�?��?Ls,��ú��׿69�]{�5i�U񯫂t�P�p��2��~66��1�%&�D`f���e
g�d�]�2j��L�Q��=�U������z��ƩOx��M�f(d�qLO��O�l���N��h��O����B�Ii��m0Jp�xZ��3��(26		(�-|�j�@�p�����K"�t��y�D�5F+(��$�pm%t<� 69&y��.D3��LD�Oc�9ǀG棥M�b"re�����;�;j�c7�t�;�����[����xn" �|J#�&B�7cvs�����~ɦ�IV:�rŶ��Icb�k�';��:���ǌ}��8V�7�ގ1����	�<��>�A���3NDH�F~��p`g���"�c�V�1}�Z��t�,|	��m���3^��%��?�&��!M���D����b�s�g��ϲ�Dx�o�8��χc��K��ۂ���0~��v�*�g/���"��|��v�_i-�3'�$�~����a�h��R"�*���T�m�yot��E��
�vgۃe�����6�[J����J]k��on�n����~fH1�^�["L�E\S~�>L�]�h�1�Q@�$�;�1?�G(�m��&Jb�8y�P�(2�i��.]��;���t����-~/|�π�V� �-�	f�� �� >xk�9�yO��Ku�v�'��ކ�۬�R�k�/�P&�a���l�:��*pg�A8�W�_��7Kmd]M��#�G�ҏ�����m�Ip�~�k�MG�ž��ȅ�1�,4^.���e*��$1�H#����N�+�&���K>ٌs��q�I+�u�l��M<J��|��>"�N��%��4���+�!HL9^���g���ҽX�׀<R I�Cv�ћ��& ɗ�onZ�6�zU��IN�*�W�l��9ۖ@��_A(�~��U�y�\���	
�6I�2����h�1�Uz�FZT���wn�mkw� �:Vn��V1��e�<���� Mru5�)����-{�Ȳ�"ǉ��m3���$������Mc`&B�0Ζ�u��yA���v��3�ݻ���E?�N�C`&!oh��]b&��[����t0���~Y���v���prYjO.m#�W_��x���6;�8do�� I��;˒i�Y�6�dU�����5$�~%�"[���SB�+�����8 ο�d����X�\�����Q'���������)�g���x���9�5�z=��:eCMVX�V��N���:��3p2�|�]q�_�b���+����/"��D�:�����gJ|�dL?Rl �0���ej�<9-��H)̛����v�D� ��&g����2�fIPZ�؊y��ɼM��&�R�מ��?JE��dkh�A�Ӏ�9��ʱ��[` ��u]6���^�W����8�T�U���Q̮&Jyjj2/�H���Lل� �Iq$�&=�6�Ïc�3v@HP����d�*H�"2t^==$��t�Y�mV�T�栎(�����u��KJ+���r��g������!��_�}otA��X���6��gϞ8xd����~��A�x�����X�L�t����d\-��� �p{�����A���ؔ�3M�zgb6��<I)<�<�$���qʆ�}7ɭp�\!��z��1Ʃ�6�Ҋ��n\y���]s�λ06���0/��}��Px���$^���8�y`�lq�@��� Y��n��[���X�$�'�N>�'����)�)�C(���-A0�����|�}q����V���FI��BE��AJχ���$��Z8{MQsf���9�i Y�7Ď��!N~�˩�2��w;�ݐh8 ��
\mr*S��F���d?��o*{���H_+*$��S҈q��ڗ2d��bU�ӵ�m���5����'����r��3��P�kG��s(�N�d�!����.9A��)&I�L �t�c����?�c�q�^|n(������ݘ$�{��O����tö	���4�[�0ފ{'xo����-�SOd:���eS�H��2�VjQ܋���e.6s�=d-�Z�K9h*+N�C�I���"��}=1
{[^��x���gط-�S���Ŭfߴf�Z9D����-�s�a��F����3�튈q�����^���_!�Ѧ�H����wߞy���K~��q��(q���%�a�:E��:��P�5���Ч����˹�z@��,5J�ɭcŔ���!Q�v�b$f��)Q�����V\o_�~�y1] DC�yq�:z��m?�y�^�F[u�=��H�%�cR#!U����!��xq�K��6Q�V��7RSFZ�L�&�>ݔ����M}<�"e�%M/i��y*$p6r[��~���za�a�d+_��=1y��18qE������$@���*Z�����\�L@Xz�2W��In����i��w/Ѹ��xr��y6�x]��9tU� `Q!��G�)y)ە�����@�/���ơ��Oʺ�(�����M8�<~spj��&��Dθ��5@�L$,��r�d��������>���w�L��=���N��ql3b�F���p�ش�T:���@���Dp)w��#ަ����bcx�|�R�����h �i���,!�-'s8�d�AoDWQ};|��Xzvz%���/[y�d�n�];O^O��a�ϻpc���O!�đ���ܧ��e����ZFy�	b�fx���/�G<��h��r�T���]�+����������T�E�$���WF|���w�6'��:4����w#��=WP��0�!EdkB��pE/~��{��ӺvG����c+�(Bk?�����8727D^Үs���� �zL� `q3�H�b|��=K-!�]\$ ��P����C�A_UI�w�|!�S'jp�,����|㽤�m��5����*Q���љ�G�Tpos��Id�J��K�eg�䣲,g�$vQ�������q�(N'��OC�J&��]���Dz~�P�,����M�z�cO*oX�!�`�6 <zp����s�����i��3��`6߈%d���~;���<�w����RA>��BA���w�H�������FS�G,��\���^�>�PM��
i9��sӣ��d�6;;+�� ���&g&�N�6Ļ������a�eÈ��Rwल��=]�J�̔=�"��<��9ʡ�t^�U�>��5��u�#A@�G��B�4��;�V�3d�@"m��3��#-���Wg�~�e����PV@�f�����[(����Y8�5�կ(I�<��j*���h�ҏ�z�K���#��ċ���]�6K_�����X����>7�Ju�n4���q�.K���󷑯���7)tN e}�.w,"����z*�	��������w�񋈆M�&�Z�H60�;r�G�q?�����L���l�k�崛������y�D唰��t�S8H��z閍I�7'e��F:�:�p?:.�Wgc�.�G�P%����4����i����������s��QXg�40��YsX��IVfX�kō��QGi`��[��~'v^�a�>�X�Pg&�%(�U��������{³᳆��!�}�����i���M���mj��@۞8tç�����D�c��nRp[�����A���O:/6<�p'1\?S��|���*��ț<@��Κ|��c�o���DQ�y�6?g��aga�$s ��fjg�,(�#�6�,�	����ɨ".�_/MAHa;U��Z߬˅�x�E,���s���yO�q@@%������N0������
+V�0G�Ǵp8�*�
����c�F��|�^p���jU�V3���
%B��ӓX�H��[W��D�Z+�ŇP���Y��]�
P��m�����r�d��8��T�Oפ!�ք^���ɳg�'EO82��z�gO���⫥!�3�X7@�7�󈁖�h G`$S��W��/n�KJ�v�x�NҜ37A,�8����7�@"&r}�("�c�~���r���]��6I_˞MݱK'n��|�{���x9����lI�?LL|����Y0����%�i�a,�H$d�|�ox�p��_��#��Fw�f�`0(F�~��_�'�}��}y{�BLN�,���`a'��q�G<�ϽI���ģbۄE�o��}��Z�N�kE}w�[/�s�<��(���ι ��[�k�Jn��G������j��Q=|#���X[���D�q�,�°�Sǅ���/�u�9�A`�'���+��zf�U?K.1 A�#�8���u uK|��8���%�L�Nָ�9�ɢ� Q��Ҙݜ�.2Ω��)��3N�6�Q����fm,F�zb��V9%Xj���͠�ꢀ��X�w������<�Ќ�)�<���*@Hj�m|�z�\?�-�F.ϓ�R?$�A�@ڔ��~���ֶR��GI�w��P>�J;3қ�KB������~,��)�EO	�c H�'n��C(��0{���ajb.��4ɏ�]x�"r5VG��ߊå3S�(XѼa:��Y�2]�����O*04�����|��]��̜'I����,~�DT��ptҷ��)��]����� vu�V����w��"��=qw��.�"�6˞w$�El	=r<?��%8�c��%&>��Tm�v��
��O��=1�W��mWF_y�T� �s����S��Oa��́0�'���cߗ�ş��.|�`S�S�bؕ� .�x|Ό];�^Nޅj�ZE�%�޽ �@���~$��y��)r���iD%�%Y��)��Lt1	���EV�|ku�v>Ͼ��oFYX�B߇0��(o��x��ߋ���Q�"zP�5{~,�ƽ=7fL�n�����eVk�+-���75�E�@8���֢��sC����VB�#�m�7@�I�j� !�*D���B�H��#����L������;�Q�s#�_�xy�L�R�Q�=��@�8T��R����
��e��k%M=���@�a��q��Q}�d�@l����hA�nAMVOF��a��D��us����F��&�"��J̳	�p��v�?�O�z b(�!�WDT�u��>�O{�s[z$m��a%�K^�p��.��n��ԖM�I{����YnG��=Y�Z�=�A��D�f�p����\ڄ�T7H�Ky�%MH�gEz�󫰯yd�7��e���>2j�[���fY�)�(�Lݍ�u#���ŪZ�sZz`��LR�&���|[���]�8r1]��5�h7�9YfU=r[đb���bi2Ħ�bl���3�xӨe���	$Y�(^1#b�Hv��B[��v�J��g0�a�Bf���DL�g�g>~	�E� �(d}$HJ�K���6���<mkn����Y��N$,����Et4�V�#��y-P�g��T���o�|7��47A4vo�0�.
[�'"���Rs���`�+�n?ԩd�U��V��#v�be!�bE�h.�U��!iZ�z�M+������t�"S]UB8�R�#6��@�B	g@1��>��h�:��S��t���M1I�����S0��)@�*����b��~}=�R��{SXR;֬N����"J�RL��O�ؙ�
�%U�`{q6�9m#���*��z �'�=6�Ͱ���E;���>{Bv�迊+��x��w�<�5��Fv�VRK�6�ۜx��	�Y���?�U¶4�#���s�㲜�W�Y���= �&��}�8��-��>0���͉yQ��*c����_�m~8i
T#�^jy�����A�X�Uz��L
��� �QY,O#�	 EVV�+e�'��.� aUb��`�v�Ow�k�r�O�HNѭJ���S��" ���~r�0)r�h �i�1)Fݳ�Q񌗼�� FE��� 1*,j�����;����5�k�U�H�
�6�x�
���o�s�{n�>�!�m�P9�JrT��Oހ��
g�I�1G�j(|��{v��$��P�Y�2N�r߸�+_���:�� �X�2İ@�i)+��7|��x�k��K_N<�	%V@L(���Y��ha*���z�|"�1������V�!V�����S�����p���
�����<��ر=M?�B?-5�[�<��X�^�}zU|���@�4��T�58�:�*�������o|-����+�AR.�P5:�
�f2�n�$g"Y�0ʓ�Q{TD8����I�q��9���G���xe�Y;��c~�^Yʄca��F:p�ѥ��O�%���K�i�?K.�&B�D��+kJ��p�m��Uv+�4A W��8�W�����1;x�ؽ�1O�`���������W�=
����)����cl�'!H# 0+��'�}`}�Z��7ş��|N�Jh xe$)]�� ��|�03��~��X `X�J��NL��A�|L �NT;>�hM]���d���>�[��č8�M��v Фk}0rg\������[��Yq�~U��;��1Y:�<]�*���@T��}�9���]1vx4f&)+��~���{v�aT)"�#`!�����ؾ8r�P�H�7HF! � ���?�52��K!��X��KQ�iM��H��ء�D�ʻ�9$17�Y�i>��/�Xys4�� ѩì��{��Mʌg7"E�1�>iC�ߟܫ̓+aFc�^���N+n٫�x%Dޡ���<`��"�qu�y�__��c2�ȉSc>[p,.��`|�C��Y��"va��U ��nP�B(-�i���o;7~;�:�,P����r���t���`���ȆmJ��Bq���EOr���c�.�X�[�u�Ø��I�f�O��5�~˅ݑ{�@8��?"��� #@ܿ>�q�W1͸),|�ɂδyc��ܖS�`�%$��CPZs����B�'�%ᆍ����|[��G��1�Q����@�i��)Zo��0ؔr$�d7���r(Y�S{Y �*2{r���[2�����+{U
�q,c�dx)|�
8��*�z�a޴��C�iP�y .��ƥ���?|�����4�N��݁s�_�^.�����Y9ѝ��}YxW6�g~d��)H"��ǆS���SNg��X����E����ؼys�ڵ+�9��ַ��2//7m��ē��zꩱ}������
��Yr��Ԟ+6i�{��O�+��ϢG莮��tK��	<�>;O�I�TD״��Sb�S�`>�  @ IDAT��x�
T��!���e��e��^�h�Y�[���Al{�_7ݼ=��Ùt�}��}��U�p���͂m�YPZ��^xQ�x��mN+\Z�x��x�(g75����2soRh'�	����yiJлe"���y��'��e��s��o��g�H�C�1�	���ds�d����npha�>6�)aS�s���k�?�sv��Z�g�G�p�K�.\�E�Y �4? 	�PDw�u��x�_����D�b�b�U��7�~�v>w]�^=�0����IZG����C�d��V�ڑ���I�X� ���X��W��_���>�鱿�6� J�k��R3!��1�l�|r)���sp:X)6uo���q��� Čg�cUЯ���A�+���W#�dņhh�8Tn���ױ%"� �^o��\�H׈'0�h������zH�d�4�}��q�禐�?���Ш!�j����O>9S��mߴYW��ީ��9ʈ�H�{�N�b�Q��� �}��u��}���i��+mj��G���p�ŗ�pe2;.��$E��p��V|�ꪫx6d�g��c7�%1��9���İ����c/\��Y</�����}a��
n}���ŏ�+����?ч���MAj�M'���e@�T��Y��m{c��p���q�ƏǺ������ԧHN��R7��Ӱ�u�u�&�`|����/�VLXj3�YR��bK���Y�L�A�r�n��=��$�r��F�\0B�q������g�=��Yx�
��IZ�c��9<1�
�G|LsG4�(B�{Ftozx�=�~��JhV�CQ8E�S�;��v<z��"�0�Q��)lޱcǲ�"�y߁��n���q��G?�j�ʹ؎�D�����32�8K b��4O���in6�K&목	�p?�S��.��|zxw��f��;����헺=xK*�y�c�.m��?gp$׳Lľ=�c��aN�e�>��v�d�)��S_I}R!�N|g�fC�!a	�O��4�����yq.�4q���{m+�شs�Z�O2��.����긗���_r78�,�$.?M�o���.��ZGJ��_��g��;-��y^|kjM�b~�!k�f <=�5�0����1O��=��L�0Md�"A�Iמ�$���c��*������4L����ohE��lE���Hf{Zƌ�@�Y'ܹ�T,��)D�����h-Ɔ�#�Z\t�sb���" ;I�I.{���f�6��<��(��cn�"��)����ۈ���
:�E"��+'#��mʙdm�7��:D�T��fx<�hvΦ3-������\���3��P�tVz���J��:������3���v���v�1����v�/z�.>���/ߕ9S����|=̭�f�ro�n����r?��
a�]|W0�K��e������"��"��,� �,z�]%�H����;�a�8��a��q��O˲��t?���\��,g"��Q	=E�60 �j�%0��^��xǻ�%r�%1u�њ�*�ͷEa���L�¯ �y	8Ӗ�,�mʭ��1iyR��)*��`iQ�5�TE�~SN��eO`7�Z�Hj�f ]�@�Y���N"	�uL����b�Ț849�S�3c���x��^�`ݳ2���Ӵ���nv`�>��w T�w;�{�tA�O纥�:�'>�U�ˮ�ujLP7Dh�>ˌ%k�D�$8�=P�1�p ��_���B�o߾N�5^'��;�zfUC����k:H�!0��`�8V��מ:�=SE���3��[�܋-;ƝM���!��Q������/��]�C�H�<��x9�,�R���+�sI�P/v��!f��m5�sJ),ҳ��K�[7��Ux�w��}���.�t�n�sYb���X "�S�4����_�UiƋ~�E�e��#o�4���Fu������Per����v���C���
���Cw,���������a�!�93a�
�
�+�gBS[���׆���*7����;�֜�M���??��j5^��ϊ�8-�oڄV2q�����n��|w~��t/�2:����v~Z�}i#�����c~Όc�nv����2I������0#��-{��ضm[�*z��^�d:�n�s�b�֍Hx{[���)g���� b��6�e��E�-�܇7�I��|��FG�V��KC��5��:S�xꇏt�e��L���w��v���!�E"���\e2�V��糈�q7�a������gJDx�J 3�������9J�n��PC��B��%&��%�
E.�F]O�{k<�� �.��^���A�ۯ�]�zj��n�#ahR��&崾4��"�3�����]��~a����#�SP��u�3�xD_��C�r�;s��ڦ��#��rz4�͌��zh�����5�����p�"e�()�yt$m�;�2G�� �h��\�_��+p��?��@k�����A,��an$ Y=�&�\���o<v�c6�-?g�yf�$<�	
9uA|D�@.��|�1-��χ=��X�W��Na��$�U�v�cq(|���ږ/7~������Ŝ���y�ǎ>ށ��K�}��淉�ӽi���`D�Ib��2:�<�c�p���� 3����!;�w�߅�܀��D���~��җ����8��(�f��]y��Je,
S(�Z8#�r��x��ϋ/]G=��_�Տ�Aa�(۪py�V�.�D��zϡIi	�8�X�9����WnW��1��w��w��{[L��|t�QįAY>Q&T��"qSc����j����S�,�fӹ�b�ϊ���s_~i��5��i:�zpٞ��#	��8��1��sߞ�le�?�}�[S�*]y"��6�MBX�03���ҫ��D� ҔAs�H����#�l	M����kq�A?&B]��ip�����G��k���2�ʆ�6�A<f���w�P4`<spr�R���G�o^��$R ����1�ܠ�p�+W�ě��uiN$K��F�sN��A��p���f-����WYǊVc�6�Ѹ�?y����8;�7L��^�����<���Gū.y)�܃��dLR�J�$�ojBxf��S��?zif��/s�G5V�V*­:ۖ# ��H���;��X�p��3	�y���t�[$�6�}��36��qR6Gi�N<f(��,��<Y��k�vwގ#�8r"n�]W:�;���ͧ�/ U8�W����m7���-�����(LmG�����V~����TP?B;���ǔ�ݨ�L�S[�tӇ���Q�¡���τ���Dh��6>[�$6��)j2�.Zg�����G��1����J�L�U�w����rϻ�H��'�#`�����"��:�K�H��pE�Uk߁C����Gy���?%v�>A�n��C1��7w Ɖ�WA�RO2�����j��N����Tj �ɫW��Re�HLG���y���˓���}SmOέ�C��8�pt02�;`�Oq0r�`d}��g>�H�ۢJ�p����󌤬�K#j:�A�bO�}�J��Dƚ�L�Rb�����>[VǗ���cP���k�Gg�㐩���מ�����\�%���!���~��{���~�9՛���m�{&o��jQ�$�8��o�F����E$�0D���_┦��Yv������~1{�s&��B{Z(�Xl�<����҂�+h���[y-�HL��:��UVs�z +:d>;�s���KLn���˷C��9���r���װ=�w��@⿉�<�a1�$$���Fy�|rg�G���X[@@���XҔk� |y"~s	����T��o'��12��_o��7�!Jk�#�ω����?�]���0�P�M��W�Z�хM �y<3N�}�@F����13�����(�߸����V�g��=%v��Z��a뛻��k�9=��!��t��~�v!T|AA(����'���.�����c~�g��q �����/%;�?�8޸�i���7��#P٫v��+�#�6$���$����5vƓd��x��"f.���0�r\��Sg11x�|(�rU��s��$�`ӕ��9��{�Y{,�bl8.1i�zi��=rx����-N?�q!$BGCW*���X����e/�S�/�V�P�<����'rϐ(��$MK�k���1EI�V#$ gI $��lݑ�#N)�,nK��@3^r.[l��wbrF�U������̒��X��X�{��ǟU��ҿ�g��x8%���p�b5=�h�� ��Kk�XXx����u���Nrf!�Xy���-�����~�?��m,^���6Wc�:rf�O;@3�F}h���E�'����J�"[��4�ohuD3���j�p�
X��#�B��<��r6�IR%��2���!r��Y��Q��;��S�r1��Ԧ"W�D7��	��A���$�{q����b}���������3.�#�$�8�ds�/>E��1�br=ɪF-��[���U��;3]X�x'�P嶙ѐ^@n�͘�e�U�'�Sh�486��f���7��O+"Z�9K�����#�[n�Ƽ9Un̦zL�+�� ��D�ֱu&LG`����$�+��guۆ�ʑ�M�T�P&�(lu��K�����HPR��|�ϵ���:��_�������	q"2`s�2~"�n9'�j"��؞XQh����	I�(��j����#�W�+N�k�š�[I9G~d�i3�V�Q/�HU������r��u�������ım`$nܾ?����ǿ��\_$P��d�&缾~y}ЮWIx��aSg��
�;HR22b:#&�WƝ�p����5Y�XRQ ��,�89w=�i�q`	��V6Z8�2�MmAI=��j����Dl��ͦ�P�S#9Q]l�W�F�yt%��}���8�������H��@\�8�汸d�a凸�s(�3"0�}�`����y�		����&Byvں����'�fz�jP븹���Żs��d�QI<�'Xw�EA����=��^���'�r�� �&���=c�D!q˖�b1��O�+To��
E~��ǰ�$��{b������sp<D����D�-��CLs�a(���9�5G����٣n�ŏl�41鰈Y,����'�&����g��W����+1H��yV�ã��_}�N�	��G������b�>��72���Z ��ͤ|����׋��9��ܻ�8�1�ǈ��}����"nI����1Cd+# ���?��N��d�݁��/��ǔ��c���I���o�P��(k����W�<�wx����9�~>~-�e��zėեO���pP��' ��{�H!����&���B��H/P��w,����W�g>��1ս:�O�Kto�g*�$X&If_�HL�h�w,ĩTc�Y���z��}ۣt���_������41!�T�*�ɵ��^%��c�~�ئ�
�zĕ&�����"��E���4��$B�����iAh+���?7���2��@0� ��ܶ?����O��h�`P���-��W�P�XJ�XB������VVlr���y�CH:�ǹt�p�[Y ���pv�N�h�{�c���5�������΄8�桘q(�lpg�%�u�u|Qi� hä),!˷&�����K��v|���#�df�u���&r�b�<�Mj�> ���|B�b�ú8u�w��B���A�4VzEie��p<F�.,7vn閞�C���*����{��h�j 6�΃=��x�*����B��U�����Ȗ6O��Og[���mZ�Hob���F�Ej�Mǚ��bՊr�Y[�%��p��I#��>V�B�����2Q�X�Ph[A��;W���
@a�bv����݌UdG��U�ݭ�B,�P4P����X��!�I�d�D1ln��b�d9��+��XC�����F�pUrmV
�X����cb
X�&�[�*�UU����;��z��2C��xZ�38MjH�d����D��-��2�Zr�i���x;��R���$�:Ǵ���3w��t&DB��w���/�;fE���?��Zj ��m=K5%.ԋ@v�>�%	1i�b��!�N#
��\+ ��D()eU(BPt�2�~n��Kd�n���Rʢq�i�FO|h�3��I�q�x�i�Ge������֩�ɯ�M�س�e�AT��`�H}��
'MT��ƃ!pB���
�>�S��^CAeA"$�w�}��P�2pg���Y�ЅE��� Q�l �%�����`ȗ� HU+J��,�pt���G�)�`���y��?/{�ٱ���Eo���#Yl�Z_Z+���	`VF(8F��:�ʠ����^9�%,O;wm�5Xgf��0�:Dm��L,7�7bI;-��m�È�sS��%�e'(��9@߇G�ЁM���*�Ƕ!8���:B5�.4�+��Ή��H��o|���,s��o�o!�3���o�S��p���N?������=;�;w�ݾi�{�c�;�{����_�	��I�>�:4�D$�p{v@	J��O
U���kV�b|�sT�H2k�y�z�L��(5c*��[�3��/{-18s��u w�v'�qìdh�[)BU9�"m�'�,̭��&�O�(�곫D$�8���T!�Z����,<P BU8o��2���췓ȣ�n��b�7��)�Wt��Z���4%S^�9���
��ǣ5�]�G�L�o��"J�*[OJ�Él�����!��(�ޒ B�/����Ã~���%���8��*��[�kΤ=88���l��%�q��D�i�1����"�6����.���g�x׽�w/��n���F���S�||���7��x�jx;�5�f����Ɠ.z.�����cb�+��*#n���G��X�nM��K^Af�U/���̂&�9B�<�O�s
��@�>8�����M/O���}S�W�y.��d���7'�W5�?�٢;|:�HG�V2x��=`�7�	@�ƪ=�	1�B�ĵ������9e>c\;�$.�Q�o�Ԗ&M��r'��r���X���&�\�!
 �ӆNc*�2����Iw�O6���u�O��BR�	�\Ù
3m�6�Z�;�Ic�Z��-�Ɗ? {,O�v�ksl�4�2`&�Ф=�tX��ȅ򌧐��)+�{��5��4�'T%��,~dQ��ugŧ��xۻ�yZ���&0�S#�M��;��7ĪV��>F�1��`f���c�I3����g�>&U�7@д��ױ�Q�9R�&�cN� �$������m�-
e�"Q�)��d}A�ka52o��XM�@��B �6q]�#����yrP���2Sn;�z�$W�r� 
ɷ�<��y�a�At -Y�t�-��x�}�Bc�4B�O�7��lxEV׉�߁_Ď�c�?�Px�ބ�`���7�"����I|Wy�T���t��S!:�u�wR�g�,���˿��:��\oK�CQ]<R���|&��Lڣ7��$���l��U)��_�9hx�� @ �'�C�<K`�V�XE+3�=L�b �<��D r���rbɂ�["[���T�K1([Q�`���}*$u�J??�qQ���K����s�X��@��T��Ԅ���FS9��0B?����J<��K�C��AB*q��e1i��lz�wC\}ͮ��7�4|	��i��" w��f�G�W�%��߉��#��]�ɠ��M^�~�<"t�w�}�#�5e��PG�B̫%�0���Y��d���  �A���MD��WR���tB�w��{D�&D�SbC�M"�p������`B\���y��R�s�"s����t��#GˑD�G��������	~�w�y&�ʐVb�(@T�/Z:�����V-N���G��M9f)y��0�#E#��ޖ��r��Z�8;o/�a��2Gɛf�{�v�D$TW��	��qt��$x`�ݹ'˦�D�B���Ԃ�<��=7���i.t�%$�����Ps��3,��]%H���"Q�ކ"�R�´��	�$&z�e]5Ed{��0C��L� /�g����K��'[�a�{�B4��2����t��Wt8����A���Y�x����Di���s����,��5L�L?�,Q��^�V)^��b��!���̣ҵ���~4�� �jзk��1��^p��"9�k���{ҁl:�wu7��w)�k�ӆ���1aܜ˄��m@�ĩ�Y��}&�O��+���.���{-��t�]/��s�l�x^���3��W�(�����g�^/��$�Ղ�Y�m�gЗ`��]�x�[��s���^�q�w��:���.m�:�=�+���:{���79:[+a�l�g�qT]�����0�|슯�;#��;l\do�x�1��_�CH<�~��[�c��$�a8;[�c��2�$�0 в�N��3O�I��V�в��ѬJ 8�pbrp�$ՃR�#S�W��� �p}�rhci0A�������q�l�'�e�N�@� �7�{�'E!~f�gS�cZ�9Ru��&b��,�|[�}�9Mu�����,Qd�g+�m��`7�k���������,=a��ok�I�H������Kg2�ڦI��	�h%�4������p�����=niҝ�΁��]��B:!�e����%5�
K79 ��%�:�t�R�._�ȹ(d� �ɲ�9w�3��6��q)�󨱟����	|'$�����pE+|�Y� �Wqڽ�"�19"�ʳ�יNn����FR���*go�)�]{S Y`3!���A�o~8�s��39�ԕia���̺�;)�Y�(ښPq7]P��W)��!1�I	Sa�d�Ubm8��T�јlL�f��}x#Nu��ΤH��8޶&�IB~Y��
�������T�(3��X�0�c�e�Y�̶Zx��,��f�~�uC�TDB�䆌�����h�\p�ԙ���f�;c���i��Ǯb,ĉ1�x�I�lN�nƳ���H&�(&�k�d��Q�ǳG�ђ���.mXQ��LȚq���%�X܎%$�I��ͮvLo`�u,�UHD�}M�4�����ܧ�0���tib�1���SlS�`�[Xp�;	�$�I���*���Ӝ1cI��x͸�9[P�~do�_�X1��v��xꨄ��f�2�Vym��T�	b�2vO��1�C#��;�L��� �}kȿJT��xl�4�@�S������a��*э�u�J*��ՃDɒ
�)���O���`}����ݭ�zN �[���k�E? YfB-�u��(uW��q��;�#ʶ��9Bܷ������* ��5͊��	z�{��,}�جbN��%e.c�,Y���b���F�4�ˊ&��0�&9H�^ɽba#I9=ݘt>(�DWHn�++���H>E���Fr"�G�c.��������=^,�G��E�$9��!4y�/���^��=�U��S���e���h6�K�`.U6��n�c�(��÷Z�T�82_p�$LX�
=p R>6k�f��٬�~b߲ А�u�I/���Ф$*��RC=<�'!����v,��jT4�ᦰz�I� 
]X��q�Ig�~�`ą �A\��w ���§�b�do���G�9I�����7��_��ظ��� �ɡC�	7> ��S����X��E��e�r�q���ܸ���������O,��'���;�ȷ�~��K�����O.�����g�]{���x�%�m��������q�۱��;�������o]����g>*��w�w�ܺ��aq�;���7bx�*�,8\���
�jPA��%$������_H.Le�G�O$�!��$D�g�:	���ߌ�b���͝���;���f"$��[F1;��n��o�#���\�>KP	Ǣhd��y��}�ȡ������j�z��I#xwceC�TS�|`�!���N�`��ݛ���1-�ssc��BL�U=�C�A�!Y��~�<��Z�G_%Y��6�T��b��Vm�)Ō�~,)��{�z.h�Ŧ��,G�j#���9��+`�zG�Y����t�K�1�� 	������a.��;����Ք�>w$���](+�k��l|5�N�ۣ:�5�d��5�"����c].�ߺ,�r�R7Gid-��r`#+A����6z�;�2�1���id�"�},6n�U��Em�6L��b��!q���j�Q���XS���F��͟�Z��E���d���^;Fό����r)~Tãdjc.�J�G�oY܈\�V&uBi��ƥۭ�O�T8�"����<A`���ā���`X��,�f} �k%��4u���S��!���5�.(`�p����a��]��g=Ji:��S��Z��u	��sS+g -P-+q̔�춹4����o��?&��r�X(���Iz�ӲS��T7����5�I�b�J�"ΐZe��S��Y]�,=;k��~D��j5�M���^�kޅ4�G�۔+��&7�x��6t�s��8��o���3���I�����\�����x<�m�����z��,��$�w�3!s$��k�&� �SU)�ArPl����^�/����|),�M�I��^b>�G�������%���%]�)5wG��PĜñi��N�x"���	ľ���B��cW�`i�Z�ŝ%�Պ؉2��<"��C�g��-f힙���[���_�s+7Fou{�w�����E�r���q������[c�nWv�~N����+?E�k!E�j9�K �X	!0�liU�Z�8�D;[�{�v����ݒ�S�]�s�|,u�$��) ���3d�/%s�S'���@�D8&CX f�N��v�%������j��������-���~-*�"��J	�E�lI#Rf��iѡ�j�<@윆ÛCD����Q�������g?G����7�c@dH>M�Y��203�ӻ1���u;;r�����.f �=8��aw4���/�.F}'�W��R�T�я}{�$�Ρ#c�i�G>��VҖ��4�����:���/ �`�e�����9����a̔�%�@T�[�ά����*�13D��~��ø	lf�wu��$<��0H������+� -2�8���Mٸ��Ė @F��a;kԵ˭�.�E��@�3�]�U����� `VP�Ndl@�zG*�C���Zh[bs"5O�alg��|yE����h�ٴn�@4jߊ�̪>�?�"bs(cI@�n3�X_T�}�평���v�`�18@��>,4x��W��H��3_u��g�h��A�<	�PƢ�k%��azH�8K�(�����rc򅥮�_$��>Ɗ�O�pc�|-�m�M�8��y�:�	#���sη3��]��;�r�C?��g%S?ϑ:$AG|�Y��"l��w��Tǵv7�o��D�v?|��ΐE�W5t_ꧥ)%���vV���𛅆$S��8���.��ejgp�;)�*�p~�uEEj��u^���KW��9�;��m�q���$&�f�D�c(UWo"��p��nr<���E����=a[����UV�A<3�k���>G*�rT��%Z,a}q%����f�m��Y
��R������t������&	`O�)�@�����s����µ�g�e����=꾟93���$�o����N���� f���.b_��&�Iw�!�w�f����BP�4�	g/� 'zw}F��I�K7
��� hy� 4�t ��c���б�P��wu2�Y(�����OVy�TD� D*H�ZY�NNT9����l=9>�FG�J]�X+{�L�=MH~�V��5�17>�����s,dv��{@�d���Ib�e�?/?�	�H}����S;͋L?�z@q=<� &�Y.G��Y�2X8L���ي��$�rQ»�L�CC����'s��ɝ�8ꁿ��S��	�!h��^-�O[��yݟ�q��'���T���I�y��|��d�V<�
������[�EN���l(��Eg�w2ì��f"�t�L�/�3\�G�m�=m�p:+��Lm9V!��8���8�
�Q��/,DW���I�^�s1'iw$�5+�p��4��ɸ�x��)썃��󘗇`I�x�Dk]���~R/�a1j�_��&s+x�S�+K���$f�8��<'o��T ʑ��>e��GA�:���;�3��ǿ��ڇH���^%M� B�͝X�jl��dC�^���Ć�Υ�X��C�f�P���'a�H�tf�Z�3�Io����3)����]��31G�Vc�����2��g-g��Z����e�����FHc��t�"�U��%�;�@k��K��kb���M]���(�)^ٟ������Os�'& 3�iV����V\p?��7�O��t,�z6�u��cӕV�u����ͯ��xԳ.A���-�ê��`����a��hL�dd��]�I?FB��0�T�� >���S�*"^�l��ˤ�E�\"02�H T�'3Wqщv�Y��8��BG��ǄG���g`���-���m��s��h�Ձ�J�lU��ڮ�䩵��ܗ��U>�!�����'a^_�,i��XU�$f��
8s����_�7���c���)[�B��^��^d�"D�6}����}�����o<�	���0�'�nD�E$a�F���"7����"7�XZ�3�q�G�l_*�Q�gdOn��Ȁ�Dd��~hS<J�3����KR�x����6�<�)� -�{��<ݑY���Ї�17�4`%�R?~�I?���ҏ�*��b;z�'&�t]K) X�Oފ���*T�\��Z�>Щf1�M��gu�Uߞ`X- t��l����!
r��$G$�۵dt!;\�Mt1f�'�:E0�WI�Q���ԅψA��pa�c��?�;#1����8!E���{y��j���w�6'j�qt �}BT��J"s��N6W2�85 ���t��A-�)��\򋠈V��?BQ��$B�10V����� ]b���Yn@�Dv�hH�<,]����ˌfjౄ^�Ѕ������Miʣ�,�'����Z
Ծ!�t6{�/�6aq:
GD�(�<-a霓���ɫ3��tǏ��g��{�f'�z�X�w����(٩�f=���x��H��������u�Eq����u�-1:N��A*<��� �16ǁ[�\z�N�?��1鈱�����ݣ��	D� "�@\͝:�LOnòr��`�)�6�DD�BlL�\��c�(��/�#4Ws
[9�����X��Ŗ??�*M�~��2V�n����C1��z�B �ƄIeV�YV�yģ.�c�CM�d���U��OB�f'�w!6d4$]�K(qh���_��<2}�'z�6�Ț�$���rp�;����F���`�<,w�[�����,���+�!#΀�`�X�A���W����DV���9����[E��p��J�D�Bk��BLP�B�'߄e��҂���3|�§M!����,\��c�싂���ݝ�|ץ�!#,G��ܷ���6�n��RU|�VP�ز��J8[�J��׾����>o}��Cdq�(h��0���qn��9���I��y�}�F�s�g�����?ݧ.KLE
�~A	i�XJ���]Q���:H��-э��Q<H� �(9�ӟ�H|=��3Z�� ��12'.E�2
�+J�n���N��y�4V�~���Ն�7���s|���5k��D�����9Y�����.r/V�� S��/�&���z�:	��(pˤ7l�b���!>�(y{Q�6!8�]X��kZ#�H�$nZ��/���P�(�l$ǈ�>�#}$ȆP���F��d�-��n���p�Lb==�qD�*)�K�h&A�RЋ���b��o�W�n$3�y�9��I�N?�.;�@P���ۃ���A�8�a�Pv�-�������w�OԶ�1���5ĕ&�W�r��MA�I\	��ɵ�^�3����xL#6�bo�A�$��$�ϴA�����TG`Yb�r-�5A�4 �5֌Z:��N��F�Q���Ad�1VV
���'ɬ�����}!���+ 4gD���}����.�������ѹi&�t���[W�!�_�p�޽�]b1bQ/�����]���B��- 94�X��=_��K1Q��?j.6�vf�H�;w쎫o�4֧]q�˱b5n�x���΍M��q\@!�j_���)��ptl:���s�>����?��lD���>��s�j�N�t����Zy/��xy��`�0fKܰg���B3�)��n�e��JH
|5�����"�w5��nbVL�$������g�9tD"�&j3�U �%���H��͉�W��J������-�JW�?ޱ�(e�/��#{K�M�A_���Π�E�Z&	�ph!p���B5�>I���@ʪO����Dݱ�_���N�Zsa���-=�i��/����'���[Z��4��@���^J��"��{2E0Z8�3���V�'�]��u��1a39�\�d h���a����#�b�UË�1A�(�P$<#Э'��@����0,@������l�E�w�� ���8��Bj1���q��#�@�X����b�b�*�b=gs��'d*�F��`�l1���8�5ѓa�Y�aV��p?���}8@��ɫ
��r2�g��
|>& *��E�SE,�g���R����6��I��y�C��P}��Ć�5Q�!Y��	����l�s:�{�8&h�%�[�Ƙ���`����[���"�Z\�	�5��UZ�" ��:v��<}kxQnG�#�Ѯ���F %�Pp>&m*��Aԓ`k�6ť��D^@oN�؂�95M�^�_��"����%yu��J�ca(9�>�"��ݿ,<���o�bg��{������+>��&��Ox£���=̳�>���֊�G�s��G?(윉����3(����;��K��br�.���ӽ�Qҷ��p鳋o
�e��5K`)&F�>�F���{/�-\w�ߎÙ�H������wna ��o�B��3pmg���.�%��Ky���Z����E��G��:��Ж
t z��ZO���7��H������iQ�7u fݖ-1�u,6n>+����/����=+��a���Y�y ��F$��uv/��.�"L�]룂hr�S�1�#Gbb�\ԣU<#W�tR<�̇�>톍���0Nv�u�����8}��x����������Z�ߋ�6���3�ȅe�zl6��5�h�V3�ݘ���Ž7��AX**��)xu8��)Ѫ�_�K�o}g���'E��*0�w�K��P8Ch�΄��T��!3S�!4�S4��v���JDΓyJ�E�+kʃ�d����q���ږ��}2���-G-b�4�4^���Sy�g7�{UKC��]8��b��5�z<��b5<W������v���rB}#����a*
�����0�{ʶ,1q�ŻsV���˿xe\���Д[���O Z�6���g�!%��6�IO8C��&V�A��EK��:����O~!��?�[qi�P�Qr�B>������˟�[�VN�0Ұ����99�y�����u�:�L�P�M����믊'>�1��A���hY#�TZ�Ħ�
��Y�gf��������"��ܺ�}9Nћ:^INS},lݘ����иN��i󲢏i��F�����Md@���Qk��^s�q~x�ҕ��ɑ����Oz�CR/$���Esw�\����֑����s�r���Q>s��<%�@�CT��t��`R���:�΅��U2 ��(Ff�Ȑ׋��z @�́��~l;�=���-h¹�v'�u�P�o����K�3t-d�ϣ�2v�)g���}�'�s�R|&���*	���M���
����o��;���4��ͻ������i5)b���l��'}��D��s��10�x�߇�*yI ��W��b����J�뾿-��o?]Xs6m��<�4V�x�{>�}��ػ��b��C�.6��B�ڊw��{��W|9���GD���x���~� ���_�F��g>��q��g�����s<*ſ����K����vf��j N}����{
�Vs����l\v�Ǩ���W�9�<:Z(a���o�G>vJB�i  @ IDAT׹������Ư<������}/.���c�:6S����®/|̖�>yw�Me�?��������#�SR(,S ,����HĩַjK<�/���k 4�T�
Bu0��,=l3�D!�u�>i�LD!q��U<��~'ь#
826�w2ߞ����,���ۙ'��I�����б��j}?qb��i0fh�}��܉+���$7{c��]>��ͣ�����i ����Iv��v��-g0����7x���ߋY&�ľ�S�O{Z�����O�
H�CW�z�&�ɓts�~5������.R�ᆫYS�������*܅n��k����Ȫ���	ĩ�r�.38��X�dX&���Nm�q�M9M�V`�͓2Wѧ��$8�Y�s�-���"n��G�g�`y�ǽegKԍN(G@��^*�Y����M*>Yϣ����̢05$��4%��u�S(`kSs��\-�i�I4�*�q��px~�DP-�l�yΗ���x�_�z ��\�]B�I�;���/yU<煿�`�m�}� }N*�	��/�Ub, X��,q�Jz�Tqev6=�t&�����x��J;�9P�WA�"c��O�9' 0)�"y�M]0�]����]�����N�3�]�#��}<e���H��!%�GEDL�Yv��\#���6����7�1��Ϝ.���u3��Ovsܜs�8�D��	Ŀ�ʂU(���2��'ۏ�V�.f�MX���#'��,@���g�&r�v�-=!��k�l�J(����eB�gbC�BD]Q����?g�羰�܋T�����*(��*[�d���)xI��K0ׄ�d���2r;�G���X��� �~0��T��!���<Y
��Ni���f9�R:�5(��3��|��lY�Z�W��^�Ԅ4""`�]{-��_����Qc�3�@J>��';<T@K��Bէ��RRd|n�+q�zD1�c��0��޴��^J�s��ǑD)�j�`�A'��#�fꓝ�@�'�?�.�-��"��-�Ad�n��t�:�K��q�/}��~kW���ㄻ�ɸ<��	Gy���q[z}w;;����w�k�i#qw��u�I�c� Ac�����'�}���3�x���;ӌ_��M����uC�tG�<`P�*��t��x��������[����{zj�=�+�rM�7Y�����"�+!S�S]{H`�S�o��+�gxF	�TśD���-f��s�p�1Cy�3��RD�(��U���rZ��ws��xK�0��q��l�� %�^9��T-��uǗ�t#���M���]BWJ �_#[%�W�7*�	��if+�?�
�sk��pe�sU� �4Y��
�S�+	���'�o	2�'�R�i��u��etC�~�U�:���D7V�}iK1���S�s$��{��c3�z��O{Q�WLے�/�=����X��x͒������+�j���r�ε��,T�3�e����Dd��D�$��^	�g�,�L�{�{�(i	<�'��x&f� 
1��ம7�e���e�*$�;�*)e�-��r�2ˑ�_	Ĥ?��Q��`�g�QM�w8�$^�r7� *|IRS�#ia����9�����7u���p
9�gi���}�F��"^���k�) F�MDc�b"�N`r�\���k��H6�l7��`��U%��n���C@k��haE�c��J]Y<ũ��
�Ӈ$���x���y������&�}�y��8| _�ę܂�������2�3���Y^�H�'㦷����)��Wڼ*�$��%粖;W�/����/]�i:�c�Uwj�g9V�'�8��L8(����.4?�-��lĲ��#r�u�0-mQ`�+���]1^>e��@`�	۲�D�������Oޛ ZvU������ի)U��HF�Oƀ(3���ImZ�mP��FllF�2($d s��z�t���:�V�J�K�gI�jW�w�s�>����k^Ӱ�X0�R�r� N^Ԥ#N�ՙ�R���E�$�n.m�]�J��٦*즊7!ǲF~fJ1Ж� �L$C�f�Z��{(X
�|�C]�L|�?P��d�����`V���A��3S�Hm����d� ����3ܽ3�H�R��'��'�s���{�~9�V��,4�c�I f̒�9&r�EP�A�b�Zp#$�iO�8;!jI��D(�!$�=��ʑ9��:��#� dh����At�\�[$���d��G�s4�(,m���.{4���0���������DjI�)�<E(��-U8��1�\�S9Bx��b2'W����DM�kԣ��j��0���mu(:�1*����x�,����m�%�*������K��_�Gb4��4�'��EK��I��T��+
o���Z�U-8G�Gw�I0,�&��[��Hy��j�u�>��jtqZ�5�����61"�j�`-�uT �
7:8�V�!
�	3�?@G����D��F� ^w��~�[�,��H�� �4��������9�=F�]J���-��٧c韋{���.�ϵ�$�	Y돮7&o�{π� �~�M�߲��\���~�����<�i���ګ0w�%��|IG%��e�c$p:8w�\$h���s�[H��Ƕ�^�r�h����Xw¿���IW��٘�)�+፫e	��Ċ�U�-����K3�\�Pl���kL�XB����J�P �$���2��E.�܋/~�U���V+������b�f��K�"���5:��q����!�|u����o�H��ilB��/��6��x"�y� ��Ҩ��Mk��"W���D0h�5k��b:�>lm`0'��k?�D�JV��ٽ^����K��C�L�kk��c 앲xr�����_JW���qM|чܵ	�b�Z`���uD����G�"�v��J|�/�",���2�Z�����I ՜�=������?��pG�į���R���,�i!��+~�Ո&��P��h��_e7���,��9���/nIõ�/PT!<
^g�6���S�z��;�pn-�6mj���0��C���I��D2�2�,����+���"JF}g,O&Z�@V�LUC_��Xh�������.���B�>���b�
p���H\��k1v؀P2���o.k|"���[�d��d~��3�� �\DGXA�6���\�؜�x����I�$�Ի%2sx���������OS���3@ �V&��5�R������1�Τ�%rr q��_�H�ﲙ�^�vT�S,A���t�9Cii�NP �]+F~�ъ �0�~���c�"z��Z&�#�zӡс����@z򓞛&� ����\�94�B[��	8Wb3��Dg����gDt��p������JL�Z��	���.��&a�����m��Gٝ'�i���X�ނ�M�������gg>�!%"2)�jZ�U���:��5���ϗ8{�����5SO?���=�B�-�0S뱬�[�q(�A���5{3��&6��ȏH����]�X�N���s�(�:�XD$U�.3/�6���׮ILB���ߌ2t++בh"����Ñ��Tߴ������h����SP�O�ƑO��}�e�W��k<IH�8tR���!����%E8� �{�a$��Ԯ�~P3��E?C���� �1\�o��Ո:d����wRDdIS���PP�|��C7����OL>w7:�|���}�8�!��6�L� 1+�#D�`��6��#$��Vy����Q�L��2�VC�ĸ�Jm�Hʫ .*��(��DĪ�ffh�P�#�uQ�W��)e���8>��VH,�T$�{ۯՑ4��Ŧ��g`'��D��=�u����jj�Q�|(���%8=-��o�6A1[�uO)#�V� �\���͈��op"�R,c�3\��i���.��L��Vѽ�D���~8^�{�S�����	�Yu,!��4�����DѸ���<��lİ,~��(fծ}�:-0�ө�����������+W���*㟻9��I���d���9���uD���b�Is�hn���izj:����Ba�:#�?������WRw�Z�m�}��R��G�������i��^j]R�h~ �Շ��?�Gӧ>�>��7��O@`�sg���O���S"��~�L��=D��ѭIW�4�^��_��06�]g1���<���Bfn`�"�l.m���������Ӏ`B�L�(�����kJ�����'��#�Կ���
��b ���� 0�=ݲ��:��f9�U��l�_���M��$Xy��{K͝�9\���ߛ�;�<�ԃi���n��P�g�r!��̱0QH[��{���J��MLx��jV��9��2h`�nĜ���H�v4��y��ž=�7�W�1���"}!W��rԣ�`�ޣ"„��Q�$� ����aB[ �e�t;;�r6;H���4��%�-R�B%kQ%\�Qn��/�C��T�b�����Tڝ��O%?�� �`�C%�d+�mp4�'?�e�P�����4��Qp��hi�	���r�YAq.��Ǳ(1
R!TF���y䅈X�
����PG��=X}��*�qt�=��t��;ɖ��N�U��DBY����Ǵ�!H%��{hnRK$���cc�F���a��Ů������j�X�n\G��
��]�
���wX��w2�'Eo�"��wɣ���,���s�В�6�#<\`8&���:���@.-��4K�M�3���w
|Y���ζJ*	�F((T�$\m܂bi8A5>&r�l�9�1�VQ�ДY�:�g��rto�T��W�T$+�L��3�Svq8:	C�ϖs��"����Hq���S�����+��FeC�,���.�m&����q����^!�z��)U�?+���!�e���~��Qw�k��d��g�t~�O�����L��rUGD�%��kl���p�_��U/�8��4�l��PtQ�A+C-Pŕ�8�ِg��Pb���zSڵ	����D�����-B�Wselk���?%��/�9�;B�K������^"^+L4����t�=�/�GWC��k�k��4�}�s�wZ��9�����2����W�PW���r	l�&�Ml	 ֺ�r��C[��8=N���Q�lg7A�O���p��=$"�J�����vX��N̕Jo����6�ɏ�&�$N�;\@C�=Y(K �]����D���@s��0˝(��Vd�b�A�#� �H:!Xb�D@�Gp�#��Y����c�ŚP�� �it���H{�RFA��(I�m�ϐ�
=���YtZ�xUH�I��2��V6M��`�s� "�k;6)VK�5��-��>��x�w]<%x~��ط}+���H3y�>�"W_�#��ʊ�ϼ4��o�!=�Y?����q�7�G>�DZ
��!e�����2Dr�W��# �b]fc+�3�i�f5u|��m�w�H|�>͒����@���I�1�Ȗ�1����AT�͒s��ӡ�ML��������G�;Xc��X�	�Q`��1��1����"
��5pC�� �(���l���R��'Ks�}���~�^��VH@��e5dxҾ賂�����ڛ�=�,1דȉ�1��2�j���%�T������"`D`c `7ǫ�Q�� �r Q�c��a�T�<�����_�	AӇI[NB� K������]�\^!�i-�,L�	ATGb�����BcC|�k�H��H &JY\�R�8�0sW8~ফSi'D3�ն�u����(�;�]��>�V����]��Uf�xv	�����x&7=�T�&�y�XC�U��i��[̱�;5��@�ԋ�Zv��/
��<�Ӣ�z��mMb�3�
�8����?�k�y,��<�2ma�DQ7�P*��p(#���������?��T�ӳ�wbF4�:�����N����BH"ЯGPT4����<t��PL�᭿�����SD�2v��T;r�	
���v<-P�Μ.a~}ݛ��Ӷ�Ҟ=w�O���'r��z������Ǫ�+bͨ�G6��p9x9���[�76G�y�cg\�n>���[Ł5!o���}"�;,1��o��p�V���4$���(>��[��{�"jT�BL�����A�R�Z�;pOA�WM<Y�{��E���ӡ���,DGt!s�8\UG��?���O|S1r2q|!�_�vDJqv��0�
r�Dl�2J	ͮ��ӡ��c��I�q0��$@��0l8����ץ�[H��ٽSs�`����0C�n�R�p${L�3wmM����(�����٭O�F�3�dj��V����]��O:8s}��M��8��=+��_L��GHڍ�PE��sύ�(:��{�r~!��{�Lx����D���g37T��2<�n����"pӓ�֍�g�E�1(�bs<[�U�	M�1�ӄ�8���1$������d�{P!��8�8�@^<��1i�iZ[ʂ��K�G���I����@��e�o]��LL~d4tW	���UVQmB��D'a�y �$Ty�6H�C�l�e� E}~�}�|(Il�>�/'��j�u�>�
(~u����é�P= 7��T��}�Sk����#vt���> ΋BmX��zѣ��>��$� HP��x�H���\D_�P��F˱�)�H�@c�FH����Ӡ�8�73��>�U�E9�q�x�[�R��h9V�n�_-�Z�$<�q����1�'���<&�&Ծ�F+�j�h�X�J����d����`bLT|��̒�yD$	��vꑑ��dg���F���>}�H���|�_�XG�bM�s�j�NT��6_��f痸�U�ni��~������p+���p�ys(�{��
�*����4��	"�O�|�Ө�Dĵ��0�
����;�Z��X��c�Ap&'�ҧ>�����5�$�(��Ŝ0�4��@�O��X�:����Iͳ�-�Ş;��l��!V����/�C/��� �*޶eUp�c�W'&D1u_hn��B�8-��$��thk���sn�
��TE�%(�q��ZPV�aX�!��q�8dc�$�� r�k
2<�"_`3����~�H� ���&�j�Y� 4�
3�8��P;�vS��@����Q�ϣ������c���y�&[
�ÿ�t3���<��GC�37�J�;7�q�����=)�z���YY�����F�y�{���d�!Y���������t�������O!x8'��7Ҫo�5	��P,7��M,o��jꈧ��l�(�E��D��`ɩ�[����q�t�LS��62����5�����Ll�喻�&���g�==���AfN���&���=߀A��k>���p�>�/$"��r���ވ�����["��"Y2"fZ����"9N�7Qb!zf����wg!dA��ފ��ܖFW�i�'V�iv��;����U�{"�狇p��5�I�3�ޟJ%L�=�H5�S�=���^����yA�ϣ\(�V��>�?]"}5��|ۑ�k��N�C}��(\������0��6�[=�ua[���v�qM�`�,5RE�ҡN�,�=�m�"��9a���!a����#��0�t�-U�1J�"攗�L�`bM>$�W(���>R�9���G���Ҽ!�c���[���_Z*�dM�Ob�3���g�P]��`��p7�]����BO�o�>�{���Uc�Ȇ��n�}J�5��'�Ƣ�B_�L~�kގK zF���&��s����,ea��Wގ�=�r�����o�Wa��>�ӘQ���_y*����������7�y~"��ց#)�q�$�o�4hí��
 ���m�EN�L:��˃Úɝq�����,�~�7��|�#Ǟuc9.]����ALx�@n���e�3f�`�,vwf[������;c���o�`A���@�gW9*Cq'>���._������n��1a�Թ�� ��?\�Gǜ"�2=�U�<L���]u"S� z��?����K+c��mdI hn�n�������'�ӏn=/YD,TT �ԀF�l��I�&��ׯ�"D�y }��B����eذ��A�!ڸ���#.w7�T�bh��2F���sF=�DP�S���w�	��z0{�@�纤�'��N��<w0�(�*�'D�zk�������]��J�f�0
y6�c=��nk�c$ÇϾ9q��Ϧ$C�쳓ɧ�[��/;rz�����LBo�����#R*҉��~G�1vܘ /�U�� ��hwV�Û�E�ݤ��?�=n�B{�����k�p��_7�0f3��bV5G�l���	�@�^��r�����j� ��d�S���\���_PnI1#��2���d��[��������~�ߣף�o�c<W�����%�����L��o�V�GOͶ&19q�z��č�;�9t��.�~���=��2=�b���b���Ds�!j�����]qյ�qNS��\�!�.�k�1�`�c���l~��aU����{��ގ�7>)/\����I�z����>��7;V(�@�  r+���<�Yd8~F�oQŎn��{���!�g=��c���Oٽb�t/¯E(�;o|\�ǌ��ᗂ����F��üɥ8���Ť�����>}λ�{��~/7�O����s����^�{b����tQ�`} ��}��cw}y[� �ݦ��ñ���9;�D�uk_���w�Q3t�7�C��{�'ᓋPg�'2�wk��,�$�?1�����gv���V��ځ��/U��O1�ۦ ��i�M�T�����eRl�Ol�;�=�w]�39Q�<~�O�]����y4��� |�"?%q
HSћ/X�y<��[����G�O�F�qe*ȣ�ۦ)0m�ҙ�k-����I���M�ҭ�U��{�����KBa���e3�#���.�������9:b�;J��^��M�D:N���9�[��}�������U��&�]���tq�>O���LNҧ�.[ ��l7ΈH�+e���FX�(tm���M�����>�k^���鉷���]��ŦM�Җ-$���]Ϲ���}���S2@���9^^Z�z�)�n�z��O���~��\�D?k|�����s��>��S�ș��_N���̙���*��66QDy^ ���'HCI���`C��г��z��G<"}���Ly���ŏ+�k�4}ы�Ho��_�0p�9�@�;���SE�I,��U"��0ҖӋ���1����o�9�x#b�+�ݛi�\n�?�)����r�w�	�k��"�d���2v�NM����졳Yԇ��j,�aT������>]b1W���hU�밋�A?	ó+D(�Yd���ua`TY[��`J4�f�|$�'�_Y�:i�Z\[��~���8�����������)Zå�ݚ_�=݆���"̦�g�rx���$�e���)r�bD)pV3t�x6{B:F�["���#J���{e�!��}�S���X�����ߏ6/#^��n�ZP̬��"��Q���M���d�y&ʥMd͟��KKc#�0G<K�@8B�iW:i��@����}�^D�s�go�EZA|q����rx�B'����-�a��	qJf.3��GRo��]�=�g_t�Bn�s��9p�KB�I\���9Q����m�Iǎ��)��>�������j�L��Aq�#�	Q�m�~��uf("�u�N��@4��Ň�<j10B2��Yń0.���yN8/�p����m	�J�$����;��>�l���5�����g6-):tvv B�#�p�
�<�y��z�=ñq�L�qqL�6�q��j��<��\�;�:]���խ^_�����l<)s`b��eOsd����o}12B��9891��@x���ﮫ�"<p!��5����\�~�v��9����J�$6h.xD��6b
C�c�;�-�;� /0�0u��j,��V��	�H�P�L%H�!o)M�n�T\&u{�boK�Λ0[�B]���D�/���t�O�B����b�y�O<=���m��}���>�	O�͸���d�o3�ir�R��\��^��w9D��0<4�t�xFG�����I^�c3=wF�72����5�}�� $:��ς�]��k L���d����<-�hE:JR�-v��2Tx���$�t�P��E����* N�R ��ci����~��?�t�M����ʠcp %`��͝,k< �hM�@v�!~6����y7tb�I	h�r�}Ie�Jq���}=o��#������^��b�@��0��MH�ę~v �%�6:�N8ڗqU	.h�I���&�G��9����Qe����K��1Ls�=�I�a;7�Q"����)-�̤���G��igiS�̯�Q�)��Dʊy�wP�+��~fz�{��sV!&p&-R˵�P�tG+���/N��vk����!V�����b|�ܮt��$��d?��)�X�[�Pc�L'P����n�-8�Ç��ݻw��e�VRP�v� 7���,����`� m�oe�V���Ft��xmb"�Mʽ6���f�|�����2H	2N�0e�ճ�+idӎ�Р��i�Z�%)s@�Di�ey�����'��?�	q�]@ y�;ߑ�f 8,Qԧ�dh������=ZP�Iw��Q6w��xU��2@X'dh�ܯp"56O���`�r�;���Q�9���zĢn�3d����ԃ��)hʘ���c��}�y��Z<�r���<!|��1��,!F�9� 2m�P_���e}+��uw��ޯ�I-O��Z���Mi�RU�9[�8
�-�����ݜ>�W%�	� gC8��)w	�W�Y�v��_�����N�}�������ݓ�
�ɥ&4��ɴVN�y��m�mm�*�z#�k�t�Յ��у3�U���F��$�n���E8�6b���]3�3wkL�F�u��vMb�h�O�I�9������ifq>�>'���.̷Ȯ�I�}���vi9�B�^,����Q��V3��{��OL���1A�W��]\\L��������7�78�\��=�<8�u�9� U[]	�cՑ������ܟZ��F8���%/�vRL���k�ү���ٖu� VD����-�~x�ܒ��}g�����&���AOr��,�Eb���u����>��ٷ2[�7_~�vR�
Q@�uV���|+}��>��3��h�E)�&p2���Hsݡ�?���T=�/U!&u|R����~���s���^��å�f!�D�����˟����oxCz��|]z�O���f�*~��D�&�x�2ѻ���H�m��<t��i�q��Y4�_�ۘ#^�{U$��Rw�H�\�|�#���r���t$�b���Ӡ�IL��T?_"颥���?��Tiܑ�k��M(�d��|s �1����KW^����y���G��� ����P��p[XX`z�;��U�56KO��}� e,�ĝ$-��3���&�ky���B:k�`��_zu��.u�nI��[<s��J�{�|Kz������Ҿ�|zދ��+�Hy"QwΥA�d��@8���aG��|��%"�)s�V�h2dテ�$�2ѯ�i�\��I['F�<"� H�U\����0vw�`�����9t9�W�T� _9���7���2�@-�,�'(Ej}�q��APs�¨\��++dp�0���^������B�,�U����&������<�����yAL��p���rF�CZ�8��L�J�h�� �M���Q����&a��w�y�At{�p�]ļ�1Y�`�A�[cv=�/�u:���	�����߁��\��+�Iy�$��k �tڼ�d7sTi3:` ���c
C���G?>�����"+7�3`T�®��BEXYu!}Wq	������T`q���$�q����?�~(뵠#ǾƯE�G(F���3��ci�x����1e���G�i�°�R`��0���[U�]QYQS#a�4b�
%Cɴ:4�`A$���T�6~��2�� 6���3�R%�WP
�t��SSi��6v{�%��@���tEW<���S�]#�?�*���x�M�L�Sw����V�T-��r�(����� z����4����ʱ&\g��I��rY�@�GX@��tx������.��{�[3�5V�ĝ"�I��w��"#�����eS=HEk�W��g_e��N��ln�Ҕ�C��F�����@N���$&.h�D[�"9t��Y���T0&��i�Oy2�'�z�pi93����O|X��?\��䲫
 ���\�p�G_�"�Y�`����E�����^B�I�����.��>A:(j���aW��i��AXPd/!(�����������&���k j�K&��yΟ �ꡙ# ��-��6YT^n���r� ���!����az��� ��!g�ۑ!	�X9��|b��
�k�v��T�M���3�� Av�:FZ�3��l.-�$ip1�3�l��_7�
���ma	���$��xC�^0���z�a��y\�Vl�ޙ.@0
E�\�����dE�"JltL�k�"�����K�3�r�����t�e��Ʌ�-mY�5#lj�����ll'��k����ʹ@�1�U79�H*=�Z�[��f�8�B��Q���ʵoH�ū�i���a"��Av7�cB@�TK3T�j�ꪫ�Л<�Z.}��+ӝw��N6�"1�ڱO�_r d��@��d���L���Ĝ B413Zbe �?"�X�C���H��kT�CM�ؤ<+EкG��;�$&XS�`�M�����_L/��Yd[J3Ԅ�n]%���[��'�կ���0G���Ff��F&�?~�(u)�g��S�Jj�p��lKg� ���(K��4^��hk�Z{�p������������?��T��1�$Ajj�F9_BO��7�3}��k�$k����#�G?����'=%���^������x����2�_#��2��K/�i��O�Ԍ9��$޻pA���8)Z�{���(�ʤn�e���z����Ϩ�#��5t\��1>$A�z�I�K��}��5���e5��A�QXH��/ߔ�6=/-��f 4��lc�C85��\�*�= �,�KۚW�X߂ZuJN
�*t�̀��В3Q����Gzԣ�����\	!��g?�N5{NV��/�9rJp#��5�jޥ�$�X �yO��/�Rv�E�
uq��a�ˣ��^�.�0��a�P@3Ĝ7��E�=�K(���@Q&��J}6]��O�{����[a~���N���t&��D��U_N{_�?��:;"���q8���@��.|�@�C�ү��/cq{�_���{�x��Fē���L��V�W��WA�k8ţs¿�y���1%�+��D�����>��/ı���������Z�6+�p�����淼-�x��(__�ω���T���Wn)����
m�=�l`8 �<6�\c8<8����BgTB�b-�FJX�
�hY��7J_&&��BE�Jx:�5���"��+�^��,+��M�c$|vʨ�aQ�Iw���iy����-v3T�A@,�=8�CTb*�fzz*����>��Ob
ֿ!��R֝I���i���b� 
�fuJ�,��g�:]�
 ,jUL�(1K�1��,�[9J�6(>���`��7�4K�٥!X{������[P�"ƴ�pnFɌNwe5��������׷D�6b�q-++���~��w�A��۷o=n�7�7�D����E|�b��-����Bn8���Mv�����o\�~��?��?�rBQ��h�e��Yx���>']��%/y���� ����ia�5i���
"6Dm'�#ǘ�D� qΡ��qx����!�V�����Z��E���Z���:�-��M۶Y,=�ƆXCM�>�����5�Ů	���a������~_��8�}p�����t�7��©��Gإ���T�)���>p�@:@+^����v0Xe���P�F@Y��A4�
�م�⨤eG+��et��]���I��� ��. X]�F͘��t:��+i)�	�ÑO���t��9���lڽ�:4��N���I�v�1j�̌@$��N��"bSnfJ��b���ge�5D˚�ư��Y�X� ���W�����0�/B�>�J3� ���qD��q	�c��D�h�Ǉ����g�%(~��]f ��P �ƽ�AR�E��l���H�c�-鱏�~.� �g��j&5���{��}�]�ci� �\51�#S�it�^i���cbg�q�A���l6��0*�]8����%ҍΠF��gx��p���(ۧ���g�넜&m]bb*�6쨲���BaK�ħ>M�㯥�0�fѼQ?W��<	������k8]t����?�i���wA��+ V%��@���.���;��g��v������U��3g���OW^���D��.��.�0���[/{�+��CC�[{$vL���IK�b��z�]�99��<��"z���p"�7릆��:T��7M��л��j�"�g`E�G�"�x�jb��UMi|l�q�5:�C�q��>��S�� ���j�ߣ��S��Ȣ�h�cT�V��H��P!pa��o:�ù�l�
�ƸA��-����2��ٗ�KxQ�շ�[X\��b�ec
X���-|򠼄_�/��BWz����-u8�}n����t�T#}߮q��mMb���<�j�Ԓ��{ߛ��_b�X$ ��(oa��$�A��N��Ϧ�c��,�.�3 �]���B�	�;�Ms��2H���?���ko�)���JDJh�G$|��8�&��m;.NO{�kҶ�/JG��L� RŪiU�d��������া#�� zz�)t��@�]Ɗ�UF����mC@LT�dl��]D��P� ��	�Tp�۫��� =b��W$5>��^W�`V��nZ�,�^���+�U�H��8W�'`n��j�nq[���x�'nH�O�O���8��e	��t�>�M.+������]�-z-BJ������Ӣ�IL|�ؽpS�|���cW����G=-M�:��q�JP���*�,��a'���>���;��:�q-K��w�7��S��7�f"4}ϡ��~1 g	K@Ӆ=PTe7�A�=�H��v�[ڗFƍ{�hÍ0oy��6wFE�W�
���#�H@T�8g����J��
o%�@sw	J|����b'��@��%^����p�XED�ҳ���R���}=�?��C�:�{Z�f$�fgKC��
��EI�Z�����,b88��mL�`BQ-�QA�������8���1���b\��
y꒠��D��CȻl!.��yg9A�2�>\��t]��Ô��y <=�	@>�����Y������9�\�w����I":�eC�PX
���PM��)�^�N��;2�u�S̥@�"����QL|�|$��錀۷��a$}Ԕ���k�r��w�� 7�
�y]�䂢���k����xb��ŭ����Q���/g��c�&嬌0���T@4!)��Zs���-�8�����c�$�Z��a�»~7�̑5�I����,Xˁ�8Rn<-,-bΧm[v���.gİ�8&�ѕE����"�X獦�p���Œ�2sx��y X7��O��15g#� � \��z��
kv�\��ڕ!�˶n�m�뵆�r=t7UTv 4��X�=]Sn�W���}{M�L��W�B @�)�\�>��w	=�{9����#q��A~�e���l��~S4��	�,�*����=f���I]�F/��&��y��â�Qm�'�e#w�p��w�P��Z�9�E�]V���>�����q�1�|s������zN���a��ގ��Z\��+%/���3@-��*��N(�����R�m�����,�.�"��&�Vg��YXy�#F)ۗى;j�q�w��!�W��� ���2��E"�s� ��a�����T���<T�@T`<��T��B4r&M�>]̣�N����;��*rx�c	M=f�&����(~��V  @ IDAT ܏�}fr��[�@^yeLER3�R �p���cq)@fĘ�M�E�C���U�!Q<�/!i�Y���p|ͶK5�^G7q�Q$�sȫ��6����b�� H򋪑_C���hY����$
p��zxą��P���>�7VG$�c��P�O�&G�+��O��~㗻�ᴠ�q�$�\��$����r�{�,ރi��<�G&3��	�ox��� }A�?���ȝm�)�3��6�ؘ'X]#e���03OO���n'�́u�I�Y9�p /ɳX�nc�Q�5��Wu�A
,n�ݴ��&	rJh��w"����d���7����aS8C�3w��.���������(��V�@0��,�@�Q�N�7�D$�0NV)7����v��q���lK��nb�/�SQ���4���ϟH�y��\��ԥ1pq팭ę[���l��,T�n$Fd ��.q,;��<�B
�f v��7���\�G����o��w��P��}dȉ���lB���43;�)e'�@0\��Dp��%)fP��sScx�o�v�k l�Dm6����%�]�t$���Z�� ��1��v����M=X��D��R{�t'�]B)b�"�H#��#�y��t���Z<�������`)�m|�;�}�,�U�C��_v�+����R����?[��l!�AL�δ��3!8z�{��� 1R�^��:��};J�
�mO`�����%&u8����B�ݣ��M��EE��d2Yj6mL�Lj�?�!C$�i�&��Nù�+��^Hgl���g=㇈�83]t�%t�5�on���g���g<�� V��va�[�SYL���� @����,ܺ	�d��t�צ=wܘJx)^qœӁ�i��N.���H��OG��?�T)m^�B|(��/}1�	_���Mg]xq���z�be!}�_�����س��ٓ��)���>ve��5���C������=��a-�8��:��GH���[�.}r4���g�.��w2�����V5�.��طH��Ӂ �^$==K\��BI�'$�--K|ʈ���Y��]�'��Q"��cͫ�d�د�}�l(PpH>�W�n�~B��(�%�<���9�Xv���e��2Ȼ�#��G�4�]���j p(����y�%aO\��`,f,��V�x��N�v�'�kb���2�	��91�¼�u/e'�TX���Q��NdK31om�g?�	���U�5:s�dQ&G7��(����������`��w�*��������sQjO�+��oNK��H�s�X!�x��ӟ��x�Ę��1�7-����_��t�6��&է�#K���4fV��霝Ci��7����xF�gw�p��]���צ�o��C_�G��E�߹k/̅TY�&��}Q�\W'�~�x1�t�7x,|c��U캷f�RpFHa����滛B=���n����$��ir����A<�86���w����|��Y�����IHz\I���G���k�&^�gVqBd��#n�w8�x�H΂�z�8EX�<������-L�=D�ȅ��j��92�"{��8���(��f��U�Dq4�,v���������n�����
�S��r�1Ua���B�G��\^{�{��Ù ��E)K���~���!ޒ>x5I��Y\�s8�	��h@�+Gv����g�����=�M6�>��E��׼�d�: ��)�LUӕߘEά&�Y����o�1�;���t��)}}b��D��g_�b���Z�:�&����C�h|��J?����1����Cj�,��^��T>+�WFғ��H�
�[�6�pӍ��oB�XHO~�#��4����婺�1����g���D�V��H��~Xz�%��;?�^h(}�+�!U�3RH?p�Cҟ��3iLh�[D1���M��,H��#��t�7�c+��0?���R�Xw��\�:xcz��(}��_����˲8{��<�~,�ǙpV�#	�W!b5 ����[�Kֱ������GX�8ܿ��Obw��ω��ؘ��臼�S�:�.lm�2�GpfBk�qHD$4�bh�xf����Ћ�����G\�Uc�c�к��d#-�w�+����pբ*��>�)Z����i�.Rߘ��I>�1s����$&�s�[� e���w������9;�B��5��aWewd�
C�!��D;�����O�w���؉]\�3�*�ѡ��b�VH.�8�곥��	4cw}��p.	{q::tp:]w��R�/���p]�r�u�����z��<�-�	 �`(O��뾹akO���G��D�^�Mc�Y^�"�پ�G�3uh�>�&�tN~�{g%m'8nˮ�Œ�������F��W!~�=�B�/+;�#����U�D2P�.�!�@�����A�Al;�}7�C�e�E��Q�1OGw��tх�H�l�H����>B<��V��{p�pRw�	T|I���a�x����x!�ڼ~5H�ԬF��\�����Tz+z�~.A�53�g�����oxd<�Qb���^�q�C��)��8�Lµ���R�B�������/=pc��%���^$
ɢ@ڂR���uR:n�i�ҙ�ɦ�؜R�J��&��|�qu6���
|�Pْj�s70����Րsܨ�Z���%X��ᴯ��0���ǎ�2#�����c=A�٫2���<�ؽ�Dǝ�>�	��}�|��c]fQ�l���T�׈�I�[6�	|'���,H�e���=�0����ʾ�y�c�F�����z3V�ibRHe���Ld��>獐�m�?�G�CaLf��<��.o�dM<w���tFӊ��sV>۴�L��f�;�����Dm~6�%��)<�%�t�N�{�Yi�Y�2*;-'䘀<;YbRLס���t䎫��[�������� \�k�~�0y�YF2�Q�&�Ev���ͽ4����F�D��ޭ]�t�Nq-Ĉ3�Sr��M��{� fh�c7�:>���d���c��$`�[��"���#wp��P���Q`�=�Q8+�K�ޜ��X�^!�%��S���1	7�ч�����j�f�a��������'#Qu�G@-�V�{!�	E��y�2����R�QV�{�~\���Xu�@�a�0 ���C�{e{D"��K?�S�R��`�Z�)�:����!`a���|U��Ќ��.��-;ӏ\�x���������!��Y�K�t������-�4�E��h��Y�g>��A���M˷��֍�y!
���#�w���gD7�Fj��hf,%�����}:��OJ��;R���p 	D,�rz��^Qi���kӍ(�[Xo���LW��i�;����or��ںc���a�Y�k@4
�������TM�ps�:"l`�#N�($�¨Ȯ����\M{u��n�n&��2�@U����D�$$=b"W��w�I ��}���	LQ��gf��$*���W�HD�<�.	.���{f��#utlS��G>��I�57�A!�A�,�a�Zn��L�u�צ+^���%�R�@�Ub�k.OW���ܑ�[��qbSk�d"J����"y�Qvf<V��v��#�M�s���[�n�8��W"<H;�ei���W������	��D��z=�1�r�!f����#��#h�z&`�2i�� r�	��p���37�il�,v��2���$��� �`ɱ@���a��ڤ4[� ls�8����ƂQh��`�Q����d�6��N_u����g�t������wn0i�r�T�����%I@��,�Γu��s�-���LQ��D8�,����!�����> r���_�|>��4����kN�����u0����1?��)Bd�sק�΀��?�9���ؕ�9Ž������ޯ��5�DB���K�:}5bL��Ǚ�z-B��������ގ�L?B/Sΐ�i"�^A�f�Y���y�����ZK���?�9��*6%9�n��\��������G�W��p5Zڂr��v�J���U��I!X�۽ݷ݄��-�W�kb9"�*p����<�x�@.�O��<�h~�	�G �����S���D��K>ю��ȡ���s�s.�D�'��i&"?I3 ��@�R�ܝ�H�7F�ƒ��L��F��"\�@�0��!�,\;�!��R
α�։E!)�A`�1��z�Lf��<�Eє7f��p������
Y��,T���r8����"�~�hN��u\�p�ru��HI()��!l�<w<V�0+i��܌��&�fL�݂�����¥� Ƽ�q��0�\T4�"Duf�k�K`S�N�J�S'?D�4�%�ܜ�/��¹sm�t9�k���OҤv�b}w�r��io�#i�F���b@��"��w���{���4;A2�� $���#�g�z�U^�1Kl�^�*JAB AhX�0[{��a&������ �.KW5���c������(⊘��e��s{�68�5�Ԑ�!�3��0~u$���-ǻ�o�N���p|h��(9K��X1��?�'b�V��^>�Lǵ�l9g%��6�\��À�g��7���r/�!�L�"&5�.�KR���O�և�L��<��|��L�W�fO��g���(��.�a��ċ	�[�J�G�0�����8Dr�����c���A�n=����C찧��&ɓ3/D>���%��3���F��d�Lܛ���ln���\�n� �;@(�R �pQ� 0�8������@ ea���3���m�	^	�."֮�dY�|p%��&Z3��6�2~�
�pX��m6��ը�<V$Gb@5b�Ӭ�L���Q��e���JO$��[ &�a�7�[�&i	S3cvg��Ib$N���g��Grc&}ž���G��U��auː�_<�U����1,����{�������{�X\Io
3�E����w~�y���a �������x��|�e��!����Ys�[pYB~��p��C[�3q~$&5�����������PkNG��MT�3�o���ڨ��C�*��o�� ��\g�-Y�����΁�(]M5�Z�VpH��I��H�؜�⪂�o�p�2��`1ZP�e�XS���Q���p�=_�]�c��)K�J�h�U����[i��WĐ}Y�Eo�|;BM�"^��=i��W1i��E��)Q���F��)_��k�H��\zNt/y�P*�WR����݂HC�ԡM��B������?� PdB[�G�B��ܿ'�8��6��
�f��j9�IH2��\��&��U�����.!�[+|����(�d�0y7��O���ˎ�$7��?"_��,�'�=o�]�Jp̅\+�������#���[� ZS�,��;�>>���"d���������ȿ�Q�<W�ML�� i�Ż��;�+������K���;!0��Sl��lV�x�4�T��>�y�wt�g�fz� iU�ʓ��dJO���x���Q^�P%�cp)����i��� yf!B��QX2�&�{\�)>#�.:���E����W#��j�-�X:+CZ�L�~�K�@�1���'��A4ҳ�p}��n��1&v�9&��"�=�ݏ��/�DG$r�B��4�"U��:Ywi����N���|���}T!�yʉ�x������prC�Z�S�ץ��굈u��g�a�;-؊p�rP��"YЁ���w�E�1P�^A2��w�oq
H< O>�hJH�޵��m����|	������;��޾����$"h���Z� �o�Z8Q��{��$��
 (��c1`�o�N_�7����	��(���A�ͮ\��#m���1�L�A�x&��L��+�;ښ���
�.�u��������>@⤅�
 4�;JM����%iO�L& ���db���;�@�(n����-x~v�/��U
'-���й=�(��ȃ�@`)K	�%��p���1 	K�l�EX�<�#�s��ѴT��$
2M�et��;��8��7R��kNyZ�,�]��)()?1ݢ�<���&�"���AX���yL�-�rpY��Ջ�S3�yG�cy�_}��%�:~ev�R��,����b��㵦��� �Y�;aW�_� x�'�#j�g@\��@�x�vq�4@&!�ϼ�$��s�>��	���*;����#
'���NEp/࣌U�,}�_�������o�s��T֔}���y��%>y��7�.njy��"�)�1�=[��ߢ<J�|m�1�Isi~]�6҂�1�Ĥ�P�wC^ٸ�(Kp�m֕3ì/0�&L!�؈�(��"��B�}��u��!�%θC��;�T��pR P�sȦ�ZATrvq_�p$#��e?g@�,~m�k��i}�Dj� bh�A�X{�(�Re-^k�J�*~�=0��ߒ���VČb t��~�
���!�a��Ev.���$�)���mು<l6����"�9��[�e���UN�gY\"Y �l�x�9��i*�qJ1CX����uC|�{^lu"���0+�k��o�#a�QH[��2V|�����;�ġ���+L���"���|���!�u�H�o��������MDɾ�g� Q�m�<wk��bc��{��ssr�=)0��zի�������wn������ ^Ӄ��{� �<2u(���/��^b_칍��XLP�"��}!��M���`��Zg�(֚����
#b�̇���h��k�Br�i�͘~�{JX�L"���ݵQض�.5��*�����!&N8��NWd�­]E��L��.�;>�ZXS+�{������$26;�1����q*�=�ghY�����]N��oFdB዗j�wb,��ͻk����4��H�D�Iܗw�i|7��$KRNEu�Fi�?�J,!�6� �6�Z�D/с�,��}:��wcER����p���  诹����QT�	B�+Ɖ�9�%�|f�
W���X&8��]�uN��d��;'"��C���$�
<��?{4��)�Ps���A����{��D�U�l�����l!T0���5΍�yVZo����G �1���ay��j�[u`���X�F�3
�܎��H߀�5��k_������J��D�M�.1�f�es�V��%/}1D�P���Ν�tF���;�NO>�e"��%��BD���#<=��7Ҭ�gs>Z�9�FO|:�s�n���L��k����%u֪M��m�><M���Is�:�$~w;}C��2c��O���n����L��#����9����쫎��]�g������0O�'@߆U�|Qz��(����8��gaFI���䙏J_�ơt����Ԛ��ĈE���4���o��C�/z��.Tw�ܢ�`�|!�}�< �w���j�آ���t�mib��E�xsx.D7�.�'؉���G/Jˍm�Ð�%8�����r���nI�C8(�ۤB�,���C7y":�D���h��r�J��Tw���͙tn�#pg5��qN�JW	��v� �e�vbr�Db$"k�	���0F|�V�h_٧x���HGD�lݲc�~���x����c;4w�m������@�Qy?���r'?�3�x"��R}��S�|o��0�-a����[��3�B~1]}�U�G@lq(�1U0��s�`��#X�����\0�e�$��_!�uEm��l��9�W|�5D�����4P�["�}�th��ν��Y�/�
�Hp�4-Y7��z����D?Ug��;�<��*��hU~j"[�#kB�d����ej�ތ;��ڜ^�soI�i˦���w����(�/Wk>{�ӛ��vJ0�ҟ��� t�ߑ�DG�����O��Կ�v�I�����:�7��A|�P�ny`��W�����_����͛b�[F�����kz㯼~��_�v�@�J�D�v������UbR����6Nq ��;�ۏ�ԫ�a��*1��2���g�61�;�id���B�Ɏ�c���C�;���jX�����?�i#��	���d������=Ję.z�2r:��gE�$N���ш|�4�Ǩ����XwƢ�ݵ��<t�����ңM�c�kj�Jg}X�Dܖ���s�|����J����d�sı%vN!��O��yV���F�1��s#]�����Ttk;9�E�z��xt�'�C&z*�y�,�`��V��Q�^&���*�d��g��uN�����%&e�M�(AV�� �L\�gM��2m���7Ap�7���O F)����M�Ԧ��(��*�O��c��yO�D[�x6�a�tʍЉ x �r��N�2�p=_�!k9�.yRt��AP��4>���+�h�!!oˆ
�D����V����)b�fn2w������݈��G�$��dr˓-m�2C��1�竮������bV��"6�B���I��
brZ���(���@qv\��T�q�U�3mt)-�"�7�fg���D�,0Z�]=��_��KY�Qb�y>2��������)f�$ָD��Goƙ��Zb�]�e<���q�E[����q04]�D-vk6#7$�D^�k2��B� Q�y�WB����1�;�F '*�i�>��ݘ����Y=��]U�f��bN���2���X�����[L��ǯ1��Hx�Gt"�_���&&�9� �ى��t�57q�1M���޹���Dm�D�mW�50��'�ɔZ$2�r�fltKZZ!}5����B��oF�֏R����a�u��Z��Y�*��L�ȑawDdU�\g�-�D�:��d�4�]v�D�E�{T�x����01㎟`��r(�&�� ����D9���9�T�YG)QM"���-Q��ydJ@�23���|�����:��c`ϝE�`��a~���uQd��+z(BZ�(�`�or- ��=u�36'L"Xp�{��܆/Q$�p�ϡ���S��Bǥ$^[H�%�㱨��}2�t������Ek�&Y˞-��{2n��Ł�8�3�����qyG���[�ˠ�*���Y�a.oA	�e� �xj��F��G�w�Uo��q��<n��s8+���1a���<c-���
c��Ǜ��S��:ĄǍ�qJ� �@�&�L��ޛ:e\��{S�[	�'5������`[Y�8����<����t���A�m-ber {-z�8 YqJEX����2���)���r���*����A�;m�}�,�q*����[i�{� �0��܉&J�?��-G��*�z���P����ȏ�B�G�"J�&NoQ�F����<�����]77���MI�8�3�5d�3�s�X�h���&�*a�Č&se�3u�,ٚϖP0p1
�.WaY��y�R$Z*v%lWY��%��_XG�_I��vָ�CD��x8C>BKR�]Va�78�HoY�0��A��=��{3�qpo��� ��PAxDK�J��7S*8�"��C�Z�CR*y�Z�sm��H�����,1�Y[x��������t�+��37��)E�&�m���	�}�cWr���
G�
����t?s�͉�|�3���9 ?�j����������o_���3��N+���f�p!e�v�"b�!��\�g�P����B�����tWdauh(a�����m8��C��� 5�4���pN%_���_%�Dy��B�Ar4��S�3���(4[H�����6ǵ��"ϱ6"�dg���_�^hCT���;�!ZUF9+��� X6_�K�|�o�&H� ����Ѫ�L�J�/��L�Җ7� �%B��SQ��j��#�JH3~(��~ͳ@@� 5�Z�Q"�%�lx��X�G�A�BNq�9m'�#C��@�}����d~%�Sˎ.�h �u��u�B*��r�A����N�:>8�_՛�7��g��Y�6Mĉmn�!׌��dpLe��ө�OL �>{1QA$$Ys�<�����b[N�R��gP^��s4XXw/~	����k�K�����x��C� ң��G�E$tt����[��(gK�8OJ� >��rO�Hu2������ ��d���1���	�s��.8'=�������� ����#�Ո�7����t��!�-�7�ǳ1V�KX ��uV�����W��Y��b{����$�`h }��_�DM�KM֊I�;c4�7��pdql4��>�.�x7�?%�n�1?s0�yJ� "2�D��~�oIv]Mf�(�����!��0�A����'?:t�9a�ҟ���b{/^��S,���� 6��0J������O�s���
D{,���.����Ղ8��mS]��nB$:XϮ����Mߺ�uc�p���!sA�Yp��gdV�u�����>�w��h����.X󇀻��@��,1����5/<�bd�����r{��][oA�?g/'9�����@6':�a��Yt����]�� V��Y}F�9J� qk�F�(0�" +A�n�g�:��݁�A�;??wܳT��n�υ�y�b(����Z��Ł���Ko�埦���x]�#�
\R��2�5UG�M�˕��<*]�#��c�Pg�?���ܳG��y+NYs�Q~c&�&\�bfr&v�2
�Ap��.������} �Q ˝����p�sJ��0��s����x\�D�e������X¹S38\aƬ�oK�>���?~��XCƙ�ME-�FQ��b���_xy���d���e�T���]�<��q�Jtw<4��>7�DDr�u	P�������'Ӄ/��x�7�����+�@�y
����ܝ����m��}���2RV�b�)�����+�	W�-Q�ě�=�;���x�[�o�~����WV�6�:NY����,���r��8a�8�K��]��f4 t	��5X�,�Lʐ��
�l��<�w	y�~3@��w�#�D�|\Q���O��,��5�fub2rut��.�#���}�`�i�԰"Q]�204T'��9Fx�$��N��mDR�;�OM���/����&��쑽xB�?�W��'�o��E���"���3���O}�����+�s�k(���v��5M��1�����O�Hx�����?;]�ϝ��!t;�F�����?��K��7ɹq#�K��<?��BJ�Pi'�Q���¡��Q}l�PT
��Z�&K���z���/{��4��㤼��S=��t���0cT�!�ߞ�����|�3�5:���
��\2�Z��"D��$���:�N��@�� ��RmS�	��q~��_���xeZ`C��\3j%���F�1n�&�F��-*S8s�	j��I�)p�ů�w?��{��n�X4e�!���P8�"* ��v{'V0�W d�$~q�d�[���7�2&n���}�,�IH� ʠ:9��ɭ��)~�w!�5?z��<J���,���=\����P(��;.G"+n�$�2�|xnr���	����G� �x�����y����"�ޤ�6�vp� c�L�����k
���rg	�y}=(�1Y�w}�bF�i�|(M��>��=�1�J׿�� �!��S�D�`�%=�@�:�z�Ǵ:���GP8��"A%�Z�����z%9i8���*��
:�/���N���}_�`Q�*]HR�l%�Wi�dTp��:8}8Uw�e���(�g�m�b��Z��ؒn�����]��e��I�f-��F�6\�3]������C��*�a�bU��"㰅�'!	�?�~�>��c����u=�r5������}���[���E�g���w�{[��t�,d6tF����+#M� Q��K %��EUiN�<;M�b�!t�2��@D�kd9����(���Էy/�f $���VI�惔�V��B��^���}�y�Y�y|>6ML²��Iby(Y*����� *������z	W�gRy�y���V�E֚���U"��s�F5��h�����r 7��۟��g���C4���`^NdT��#=�w3^Xs�d�*1�Ӫ�ei���L�Gw�e�j����SG��.���kM��ʅtƦ!�!�a�7%���2��f��jg_N��͎T���T#!S�[�mF'��s�/L�(5o�����?`/R#�]r����i����*k��4ٺ-M�f�=�o�5����	xh�j/6����c|{��K�k���{@�Ϊ��~n�wz�L2)���@� �K�"EQP������	O��O�. �!!�I�mz�s���������ܙ�I��>}{��S�����Z�[}᷋�6���"#�!�O���DW�ŧ�X���H��U�&b�#ö�!���ǲ�G ��	�\,(�c	s�B�ܢo�!�*���dn}S��W��g��2%>ՍT�p������u��̺�����'e��J�-�eS�>!��Y�d�e��.��Rlʝ���+��v|��_������J��k���G�a�w�m�|�V�y �$Y���z�� ��q�>��~(Rc/^�/zɋp���@�w�72D���Dc���z�p�_4�*���G����&g�\�)��?=щ�gb%�,�s<ăpt�g���:ۏ�u
�Ċ5/�JD�(���i\&CX�nѸ �q����Q�Y��ƺ��9�r4C�0GÝT�^�U[G��r(z�%�1��*���F�$oA���#֝F0$ܞ��2�k,H^܉:c:V�~2u���b#
�&�*��:7Γ�l��f�oi��[ӝal�@$���Fo�b���1p�3!�x
�����g��8�z�hR/�������RT��|�8��G���	���(����+̎C=c���{��}OL�e�@"��"H2˝�[����b��T`���	3-������22�զ���~�/o�|�b�w�΍��l�}"�ތW),AD(�p��HX�-z��<Sw_GսE�����dx��q�w?�vW��}�Gc���OZ�E(:��A<3ȈN�"w��E���������I�E�Ϊק9_M�#w�ۻn�N�S(6�%��ը�NW�����a�<l��#=�����"�.�9��}��g��n!&�K����+"�ꄇ��&��*�4&��2��=��(A��8�<ey[MP?�e�u0k�xf�O�M`��K!`]�l������y��p�<
�����v�r^c�LqB��S,Lcx{._B`&&�wc��#[G�qԥ=�O�_��>"i��$q��<��93��4L�[s1m3�Z���������ɘ'$�q�uZK��.RpeD4����Zw�@h]#A�K��/������<��D�b�]W���{I|tO�,bN,L�'�W+JO�s3m�#B8Ҧ���-��U��(�a��!���^JƉ;��}d<�G�K.�Ǹ�ƻ�����d7eW���Z��Y0eKi9�O�H�G��<3?�w!�	.�*Z�|��p&7��@� <~�ɷ��.`�m���~�M	�Tİ�b_�W��ޗR�x5������+�@�`�j�Z�jL��(����Ǯ[�1��DQ��z�(Ү�$"�L�q������?KN[-Q�B������G�!r�7�#^x��S*��RQx�TK�b`s��jF֞�^r[���\���@Y��4�:���<ɨr!܎I"�������E*�Bu2�Xc�y�-H(g.�8V��'�!&{��O&���{d�3�bA���>4��`��Yt��D�Y@w���@�ţg1�j�	ɳ;�A]�����]j���������������{l}�ư,��d��W�D�fd�lz��x�w���6�q%fA1�JUj�����)!9��p�3�f�v�ꗳ+�(��wq<r�Iq�ş��uk|��_�{6��sn�#�@Bf��"�ˌ�8�Y|�SJ;�� p�e����ܻ�^����!^8gL�V������݈e#��e?�rR��ᵁ.�dG�G:�Y��F��y?��RD�b�W�`����;�q��?�$�'N@�9=M1� ��9a���1�۶��$B�&���G�k]���d�[�bE졄�$VM�����t��pE��4��O�5�AOw{vc�"�1����웙$莴���1�b����ULQ��F1��jzx"}h�Й~096;�E��:�z&g�ir�0	\����߼��I-er&��p/�P��?֑��7����Q@���]��?p�j�
�mv��Շ+z�ue��=`)@^G�Z$.Ƥiga��������O?.��������.
;���	#��y	��/�y��0�^ ���1׳$Ƒ��ZcL�[E�W� K�b��}���)�UF�W��{�.�<n(~�7ߜD��'�?�i|&��4���Ϩ4!h�d�~�?��LJ���������q£V���l"�2�
��
 ������}g�[{||��_M�����gfrE'��n�����wn��xW��Q �[R=�1@/������N�O|��d�Caʜ�M�J�e��F���+���)�+�UD$+7F�Hs�́ЋI���/�[wO��z'	�� �<�%��@E�~	����[���wn�y�Ek�\7�թM��pR��Z�rQ\����6����p鑘VNxv��q���cOF�{�$�t���L���T��'����S����D���p5�/��h��{w�=`���5�[xf��w�!ϋ�ˉչ2Y1��i_��_Mk�]��߅��%��a��ܡS D��˸�`uW� 09s���S�r'��0����K���M�D������U���Sw�2�F�z#T%
U��T� �{�dF�1���Xvʳ���m��w]��X\�4h�$��Go�b@��e������gK:����A/,���[����w����%q˽� RU��R��ft��q$b"§�<��E�^�h�"��|'kN��KN�v��Aj3�7��'�4�r|���|�&<a��@�`�����F�O,J���pf�u �x��[���mv�:��=7��F����oш^rݚq��8��3����G�����/O��X��&��6"PKY����XΘ�[o�k.�(�K=x�"
���"b,�~����n���l^N?�������.�U�7
L�-U!����c������ �O&��ņ0'2�w<�Π�oe=rM]JR���������1*�	� �{�sT��c��0���������m]8�������>���ām�I���M����\t)�(1��p��4��� ����L�e
��k�9CV�4g>Ӣ��S�sP�m�'>��8�J���Q�#�O�A�7������Se�C�(kΊ�Rȕ���� ^fxݩ��qO�m��E����q�Y��|���� <�I��vCk��gq��*�::�:K� n�-vl�O?�q��&~���6n��)`Ms"���	EE��@�K�u 9�x1C@���kr7��e ����0 �#�T!�y����[�ݐ���m�h�bN��p�D(=�&k�����X��er�"�Z�f@�@6�nVw�S�顣��S>,5ʈ�&u��!L�B*�Ql�0��ɓ��]�F?SP��݉#Q^���� �!���#$�Ի�r�Xv����q)�Tk3V�Sq�A��jU�˰qƄn��iΤ�#�P�:�sX�f)-R*S-���ClS$5��<	�+jjc	JX��P��ԁ�d+��92�'}&��K�e����M�>�?]X��&�;q%�rz �MC� @��P�����C�L�̔q"�A��jt�"b��bcOZ �nw\�u�#���x�ѵ��|�Il��S������n���X�L�����`��ħI���{<p��`1|5�nq�R��
OoP6�	@�+B�6�d�i,E*����a�l���e���Ͻ��[���q�7'.IBA1��ۺ�z��-��J��9�m�T��/����o�c��_NCQ�ݐ{@�6���*)�I}8)a֬;�Y�Y�$;�	ĂI�ؖb|�h�B�)�w�j�G�U-�Qg��!JE��%�&���@VC�Q�]o  @ IDAT w�.�t�y�8n4rIE)�;�L ����� ��� !�s8�����a�~��Gϳ���胘��;��)UYZ`Rʌ�5HmX�,ͳ�b�����:�Z	A��f`��k��yz�Ns��9���� �V��
%�\���-����H������]*�ż�Z��D��A��}ǂ��~[���utl��54D�Y6P���[�O����$�	��{��
`���.X���Y�F0�-_1_������W��{�d��Ei�0�X��Dg�ZDuQ�_�8=��Vb�-ݰ�A2Ѣ_���J��|�҉cJk�=�����Y��E�};��A� ,�wP��x��|i�|�+�W��ص�}�WH�����R����&A���}y5�r�1:FE� z5d�T\!1K!�Ġi���4�,G��[�Ŷ͝�f��'b��:��3�H�Z�Gb�m�xw���v����>.��3G�4~�����ڂ(��-������K�|M�3Q$��qT����	����xF�ߌ:�饲�i�/x�4.{�
e��+m��E�;��k1�!���X�+�@?TD	U7��S��2�! ��?�p�Ca�m�I�_�y�ŝ��:_��Wc���� �m=K�`��ÀRkNY*Dog�#H��+�$&��@�Cp,����m��h�*X�R|�o��7�s,�n�%E��^�M�-ܶen�7�*(7@�t���J<K �?�`T���=Hȋ�����{�C K̪�.0Ӗ���τ�6�9�4�U���,�[@1��{�@�ƪ�g��?��xѫ�@����S�B��Z� ��"�>)􊶲�wE=��,8�ݛ�L�r�i���G��
��n��.�!��[2o�w:����*p1�T,��!Mw`^�-�jm���NfX]�>Z(ų �� Q텻����x٣����й��x�z�
���Nn�g��GŘ3��D�w�^f�S�Xx/��9��^"�z@�o�)��f��k�_P���%�g���2�C�7��X�p�+V�rQ��=qy:J��HjGx�.��"����Q8���J���3 .[�"&�A�����Xxe�UW�Wv�X������On�nr������$&"�J�" �& ���;Y��%�c��mq���-�!VW���D�6�GC����Ly��p
�i���O�VHՅ}V��Do��X{fo��>��	Vy�u�O�[B��Qj�
B���3�!\nw>WbP�9E<=��`�ȏbxu16N^��T	����%)NH`��(閸[�3�$ �;�>�9@�&fr��  �#��!��W�"��a� Pz�r�f�'�ѡ��N����E���ƛ˅�0��4�i0�����թSg��>)~�]ږ���J�EOI��x �V����YLߕ����U���e�����=�(�S���i�T��GLI��ux��kZpkM���hN�z~O�}�S�Y�i�[��&6;h�nj�4��a}seY�6D����dQ�إ<���;}h����`\�����M7/�Ov�	��DN/�����S�����agRNA$I��O9g�v��_�xtC������Ѧ<A��)��=XiƑ�����T���{H��	�I<t�n�}M����Ź�1��O�v�Z7]���x凢6v\�nD'e��:	��k�'�Ś����b���i��}(c��LkH��~�.;0���6�㊸�{��(}QF�.o��DDS_"�f��z#�!B��LqZ��?"�rs��oI�d�p}d����񱏾����T��K�[�^�o+b�f?
�w��먫�|������!4-�k^��x�9gC%�ddD��Y��R#)�$3��g?-~�e/�7t/�v喚L��.ű�f<8^����X:$�Q�H� �>H�kpBXq��_x��U�x)a�%J�Z��r��{,�כ�7��8����X���BY���Jt.��|�Y$�~:\W��9���2�PB���G雹'��I 
=�_��$�n�I�ϰ�)��6���_z�q9h3�
���z���%&")�X�Tl<!Y=>��w��WcϽ�R�Ӥ��$���z	HU=��X�ߎeO����\�t%���h('!9)�e�f�l��l��^�s7�|Sz'��o�f2�o����Nύ�����&�+Q2�\��:=�zܳc���{1�?�wd��Ĕq�	���ј������~8�ZL2�)v\�I��l3uu���T�O}��7�	�!���(W�r�Ť�'4ٕ-1�N��<P_����B�111�U�Ca^F<��gŢ~��t��[�e9�&9�A��W ��c��=�{1DF�/�}�1D�-�P4(^����g�ft08��j��ⱅ>�z�h5񝜠�7H��,�Da���f"�T�h@t^�5�x@$�pA�@�Lˡ5��.oe�&J�s^p&D��l����'5�^��7_�6�3��6�	�Ң�Y�w�R��L��Ԣ~��ߐ�7k���!W�<�N�v��O�����*�3]b�?$�!w���#�d�$CT��;멏�S����+�9�{�q eLi8��@��g�g�ǡ�X�������q.� Ȕ�,� ���8	�y]�<����T����N��CoU�&�Aw�l���-���l�ʸ�i�O�
�b�#Ύ�㞁8B!�G����]cN6;Hε�w������| {���� ��	m��:���������?��?�|���C����o� 7�����
��V�^�o0�([*y�m�<��������^���1�%��e�~�-)Ҕ̔�+�?v�[������<�$����`<3X(��Z�ri�I�G��s���8��8��A��լ�U2ĵ��:^�K��b�4qR��L�Q���e�c���x�3��Ş��-�A^ڨ+����[6^k�#���QB�c��@|�$�6k�8���qc���5�x������1(xV��L[�֕�;���>�-�Ϟ�P�C[Hמ���qG�a.R0ˆ����X��C��F���lKL,�`�@�f�<񑏊w���F}�EqLu��	��!��_W�Ga�3������i�B ���8�9��_~{�T���;u��\�D,@0�a���	N�k��]Py�9P��@@M���,��7�
 ��PE�ڻ6zOx�da�h`k+ g��Wǽ��0���D�����YA!�[�p�#�O������(�0������Ƽ'���F��̠�?��	V;��+����;Nh�&6_�y�W���c��$0O�$��2��d2�?e����XF]�t"�FN.��g�=��4*s���?g��
�Y/I�1@�q�$>'���	��ނ����xj�d�j���q~�7�5����<f�ŋ�b��'�TM��X1]�;��T�꯬���[7\�2��8_ �AgEf�^�Q��)|Z�c�ڧ�6jLw* ;)J���&��;��v!�
Z�	Nϰ������?�-��'9t%`��ļ����3� C��{��d�+ �;���'��s��c�Gg�b-v��8UA�|5�ɶ�:vj��`�g!DM��e����Q��+�N�D)	����T��X������$��,!����$�d����S�.RG�p�W`�e<0	:ĺQ�̘�P�Sb��	�S�@���D=?�r ( �C��r�&At�wA9Z�����f���⸣V���N?w?�6�W��b�o�\*�5(�&�B/��"%7r �}[���#�a>�?C�.�S�Y%'�H��[�BP�>��(̚@&g�<j̓����&� 9dq����6G{?��{=�+�TA9���D���$"V�8̷,�+���3����b�����O�*� ����%Dib��N�n5P��v�U��j c���c�Ap�Yk� C/2����z+�j/Z�R���)
�W+��m0�SԏTX�2qX%�W�jC�d�@�IOKʲ�|��k!�M�B�VD+%����18��g���Qn8˲��s���v#�eOw������s���y `3�K�=�g���{�'�\,��ý[�[�9�S�T�)�8�]�2���시n�~a�)���=��GE��/�����b�̢X���k�ߌ�G��"�]	��S�ۢ4�N�ĳCA�������3��a
�@�wy��"��z��Q%q���oI"������������%F0�vPv�I�)����`��ט�J�FQ��/��UYR|`F�8�v���<!p-�`�>���٭��k�V��o�<ȥ�I���2��*kޞEK�GV�
sq�M߈�+�W�i�s��y�%�SB����������`g%(xg]�*ű���]���b�]����^��Ȃ�2'y��(5+���4ƌ�S!z�B`��	q�u�7��h�Y4ӛ�F��Ja����� � ���z�Q¹m��8�e��p 9,�҂�u�Sǋ5���ۣ̎gfwL�U�bf-۸�IiWk�Q�XjH��`�2�"�]qQ���?$tS��&���P��!��"D�Z"�����űf��D�Q	��&ӿ#"�H�.��f%��A��(�]�/�
e;l3*���eV){��J�9�K%���o�P���L������4�)���(ٗ# ���4��p.�/���oƤ������xy��^��"ʶc��/�zޭ�����Md���Xth�����[~�NE� Ț���6������.����r �"5%��_�.�uO|~,�8yT��ɑX̎�*���eǟ��	�aB�����X��\��+���)r_ 4xoj��hN^E�>r��\t�=�B,n�. ����DD9�N�6F�}�]�Jt���>��>�Y�v�P��π�E<{��- �d<��c��@0�q��ann��L���Ȋ�M�UM1&�ܯM�5[���'@(`��n���QA�94xLL!>(F��#���ǉ��ͭ�ד�Nd�q�p.ft/�QJdu�iKN&H�Z�䡍:
�DHB��&Z�v�x�wJo�(�f��]��|+
A�!U(r!���8�(����QR��l9���f��w������������H�qϠ{b+��h�:������Z��t��sp�u�4��yd9o
`�=���z�<ց���1���K"��O� ����%��G 7U-��}ƕHLlWb皈I���[�q��'�S?�Ê�e���k��"���K�:�g^/7	��`����D�u����a��Tٜ��<�	�&&�Cg�m&w����aI�[��X� u��7�\Vb�5w���w{����y��Pr��
�*��'��6NNE��S�1tV<�g�&��Ӕ���7|?�;B�z7���;�9�Щ���1/��?8.�jt;�s�gn"R��~"J���5Oya�e=9Lo��VB��Xu�*��Lae��;�>b�6� ~i�	HG_� � ���͌�´� 9�-���ɭuoו�Y^�BU�8.�,*�=,!"�u|�3�ҧ���s�����\���d,֧F�`�pi1�A��b������yXq��0}E8;�%���Q�#�`�����8�X�|SdE�l����&��
�Pz�LA83T��H�ѠAF}EZp�=#�g'�e,
*��~� �<����-��i��4zq+�a'�!�0���^����y~l�񫤃�3���2�_-|]���J%dB������D�L���\�?wƃ�v!$:�~�:��H�r��-���mޜ�W��p�~��Pqϗj�d��$�p�~g�c�9�D?]b�@n qIpᚾ�ǂq�di�}d�\��R��ĕ��9��"ti�}�+�;��f֔{D��61�����<���ۿ�xqV(i���� 8e(��ԩ�B���Yv�j/uX��̔V�- �ʓΎ�_p  Fyh@�W��0�e���I:�.ˇ�+'g���?��-��}�}��8�)�_ ј!�S\����n��rZ�V����3�Cַ���d����1�=�ep��pXZ��ɪ�Ρ���g\~�|�[7]C`�ED![p\��ћ-�B��&
�K�e�����:�n����`,�9t���C���/},�;n�GWbǝ?�2D�SF�Q[#Ï'� ��,��K���>�m�i!a�z�K��Aq�&�Z�����/���k�{Il��8;���!��r��gA��XS�������K������R"C>�2 *��x�8��:^L���c�"q��=pC�T�Y,O�G�B
-z�/~�����֪g��i!�H@�
����x�k>^����R�=7�ō�>��+�@p���B/���๯�����l��};���3J <O3|�Hbi�K��N����X��q<�yߑ�|ӊ�8Sgֻ�z�f
����Z�D�}��r4��a��B�v���8���'�.���d��T��>Ҙ�����q����D����=�E|�;�:1�㠺^����sl��obi�6B�! -s��R��1�J�(��"�K]%��UGg��+b�3���d��~<<K�ʉ�a�dӲE��-�y?�`�8���#X�]uG���1�NGi�o��K�(={A+=C$�4*{���[�q�H�� �0�®�SZ�c;��o��}��Xُ+<��f�oA���0i�ك��0z�6���Z�7Fa�l���XSl�5��b i�J#�F莗��p�r#q3"֥�Ū�m��oE�Q������yu���f��0�b�=�/LRE�
io*j�@L݁�
P���#�Hepqܷ�X�,[gZ+��4�xQ���s���G����4�'J3p2�������l"3X��9���k	F���ƴ����K�ƮXs�Zts���)�*-l�-\�-	j�Ŏ�]�Ա��%�u���B���QbNxM��o�"&ٙԱ���n�~?�_!m�z���^��7&1�a�Y�������#�<� y!t�7�$��WC�����z����D������� 7OS0C�p�"ߴ$���7ǣ����}o�|i�S*�L�����)�ΰ.I����p@�? 7%%�1�d��POl����G� B��7�"Ƒ+u�O5W��2l�ƝGw�L�T2�>���ye���Xt�Ş��ɛ�C8"����TٹMq��xE\���$*��I���/ى?��>�����Ʈ18,/��(<[Đ� *���ID���F��<JN����E�4Q���	�f�
Ѓ�w;�!���*"�>0N���X�
ӃՁM�]8�M��W��("�ؽ�Ԕ�/X���KdT�ѝc�䅗��4c�BS�"�)	��%v�˓��25uzJ��H�#��\g��aF9���ڂ��e����p�%*t�!5����\s�0q����It��yF��X�خ�c��?1�|~��*�њS8�s�ݴ���Q私�ʢ��K(�Ǔ�9mh<�G6�O,D�.b�����>��
�c10DJ&7�-�r�,����I�5�v�W�t?�؍C<��t0�̬fPl��������� �_E��| Y�:&���8���oQd���(P-�V�t¼e��T�6�	"�籥�j{#��æ��X�����1�CaҡSs?U�I���~���
�?�fv�r�`�~p[�TD3c{��"��[b�e���M�� �yM\�ynD"b?�v�'��/�ǭ��z��ڼ@�3~�e����� ���YH���k�r��T`�U�6q����OѮ�T`���^q�h�47�*�p(�|��o`#""��J^�=ȧ9t9D�2HT��� QB$P��2k\BT�g�4��N�Nw�_��y,(.�z�f���(-ERD��A���ho�9ćFu/�vd}$P�}LGQ�k��'�wTA�Q�d�ӚTXo���`m$
~༺�8�)h:J��t��T�V��C������p�9��!<aX�T�&�1�Y����H�?�z��� (M�h�u��&���D$��ū�+_��ŉw8t��Z~�)����=�����?�w7�����}�H�z,8����sύ/}�s��K,\x�G��}u�w�h �!N�m��>���ElM �򢻼,�0l3Mg�~�ES	��vϖ�֐Py��4��aA2�F@m�Cxd���g�Q�O؉���-={�<�B$��4;��l�fp]�;�wb�5���m(������"-|���e<t�3��d=zs�z�F6o�SO<	�'�-�I���wE�v���y��@�8X��m)W��D��RY��^�Y�*��[�yV�3�x �ݣԃ�.�h3Ԭɗ!Tp�a��~B�B�,c&V���+&끋���^� L��u �fV��6/11Rw�F��6JM8�
�J�j�nŽ�]�O��wT^��A�ч���7?�f0���c�#35�i/�x�Qf� |=��
� �}H �X�6�,�EV��(@����k���D��� #6�*:�"l����j�<m�$�&�z��|߀����8��N�1�<��:���`��7>�a�w�������wI������@��� �]���ݻ�VtMJֵ�Ja8��o�Su�|�,���C����q��/x�a�I'^~�91���'��-���bR�:������~7ר�fy��i��12k�bs�����T���w�d���i�k�W��2��'ߝdB���ds9��̍��5ψ�-wE/;7ah��\�'�BҒ5�M8�Q��r��t�עǚ�'�=@<�����e!������и��M���vmЋ���4�~���e���y������s9�&�Zʨ�<�q�q��R�g��
$=}�[8qZ���!���@�2�f��Y��aW|ȩ�����"������(x��6q7bs��@=��(	�y`u�Q�h����i�,�I3����,��A'�#�l	/Ta�6>1:�e
��=�g
�a��!��}��H��r���/�9�D���ai����������s�~����j�nT,�*9|I�Ձ��e���+��'�t>,[�<�^E��W�ԡ��M/�3�
)��t�7:&�0�jݩ�ө�G�Fi�Ց̜;M�>O��ĥ�T�7�Bq4�{r
Lz-�r�ñ��t �0���d:y8�����9K�5$��i�y�,�
�]r�l/�\<�/fck1�K֞ΠȚ&��0O�o����G8y�����h���'>6+�ڜS� �'����	�� ����8��Xqٳw#\�1 s�dݷ�8�����c��i���Kb,d�
�:'`p��A?3 � �4����4:��<K$Tt%}CzϚ���+���U�
���K�DC���ׅS�Y� H�I�k47�m`N:*���^i��ǒ&�yL�M��V���}�����XBD��u����h�KF��k��k����������ݑ����y:����YF����7.���;�%m&ސ�2��%/}�����H�$�7U����?Hʼ�%j��)\'^��W��I0���:�$Ҽ���ձQ�p�k@H�l�ԯ]����C����~�D��o�����y?�Ե������E��{�����>xxf�eߺ�e��3i��b���z�vҐrY}m渚	�{�Td99ʡ�! �4�Va$�=�i(�ػ`Oa������<����'��jaJ�lm9φ�~l��sc��ɋ�P("H���7gK�z=im��P� �,�gg�~����ٻ����g�����D2){�-q<1�S�uw�lQ$$N���<�$��>x�c��{]�Lv�!�������wM�)!�K`�%X�2�y4��4���O��e$T�Gg"m��2X�.8�����x�a���y�s�+~z�R�kg"�
�^H���G�E	YS�/>6����(R �C�����@��l��4�r�9V^�_��@�D�8�pV�wEدb�T����.�O}�2����cF�)�פ`_�����w�o�,/�s?��O���q�1'�?ʾ��?�����,|�쫗��'f���&�ǩ�d��D"Er3�wxY�lW����}�	\��4�vG����z�'�s=���{wܱ�:��F�立bţ��ɒ�j�y��!a�R����?s����@t������������C�ŏ"|B�l	
�HMb<�b�P��z��٧r��kb���zwx�ɮ�����Ms��vl��|�~9x�#����k]�Xd��L6�f������sP-��s��wW�^��?�\��9��\����5��=�{|����rЈ{{I�'PǓ�*��/�*��j�j!jt-�,J���*��S�oP�%w ���>��aIq]�(� p0e,��G&7m�'���yi|������6L�6Ci]c�e��/��U\J�o`�J�p�c��΃L<$��O~�_\��,�,��ML�ɯ��1ٕ� �ʷ92�Ù b0����;)��B�BP�iY�Ɖ�z�Da'��3Ɏ���~���a�%�v.�L<�*+ǢO]��Ȥ͡�A�I�C�@�;D�N�k:��nk9z&;M�1s1����:�%���#�fH���m96����s`H  "һD��J�D^�V4�^2"���2��/�E�D�����'�p�GA�s��ZK�X�0�Z��.�֦��8���gs��?#���&|�t��i����Ѳd�}s�%����=�?�Q�Y�G������{x�~�c<�Jd_��[�^�3zw����PZJh�0qx�"|�س8yc�f'�'�[�5zz�M�h���B�������'�:���V��p�K�/�=�IӢ��B�W��Uq�7��<pA=��L�X�>,�����Y$�wb�Է�Π��R��m�S���;nY�ؤ��ѱ<���&�uX�<19SSX���k	+��.�����~9�Ȩhs��B�1J�����@��(��>����Km%���/�L���EcÝ8k� T|��:H�3��q�YCdq�ll�&!gf[�å1�VP ϶�ҋiR�]R�&��; u�mB�+N���O�}p�Sn�>w�H�ئD!��?���s��O1@Q5�q�#M�E���<gq����!�w�RvA�(A�Ö��ߧ�O��M�q���Ro��]�$����; n�`.;���5�w~�?�O4{��Ux���3�O��;���8>�%���;k׵�t�J��&�2�ǝ�y�?�����'�w7�r*N���/�����3ۨ �0�\�NS�|3�{&b�vRl��q-��à�:�.p;8��ݞ/��a|L���K]0݌�M��ՃvjJh\����>;�>�Y@�Q�ӱ�⓱>Q[�0E͹=�˙�Q!F���I�!b:A	�F��%�29 wz�{ׁ+���X��'ĎM�Nk�N��(�đn��8�̗E~щ��o3�����C,����Β#�6�(]��$"�|	ĈqĲ4A�"n�E ��,G>2!��ل� ��-��p	"`BF�c�`��#��t�A9�S�|�$�TKDq��7�N�h��X��N�7���7�.l��;�[^���5
���qZ���
��H>H|s��u�m�Ҟ�(�/�r�#��x[��{"���N=�p��LdM7�l��@��0��S6��F�[�r��t���W	�_|�I�����S-/LRB3��ܗƖ��'�W*wX%��u�鬉IrddU|]�k�r��4���s7!#��K�{}j�A�[����H�DV*y�1��7/�j��}}Q�D����G������ŋ�e�l�/��?�FZ*��]N����b������1��s������	���,�-�1=�$V{ÚY�/�m,�I�ܺ3!�Kπ�X��>�@�����&Ƈ(�
��0S���q�iG�EI�- (:dʭ�b�I�89�a0	��H�`��a �.v���p�op��':�:����ţ�h�|#�w9��V}�ȑ6N{�V������x�t\x�W�S�x?��z+��R����B8�����>� nK���]�]=v����3"�1%C&3�I��ǁOpp�w�� �.RJL��ԫ�����L���}\��V���H�co��l�toJ`U��Ν�BF͐�������?��x�I���A�J=D��zt׵�yz)�w�l.���11���F"$ݫ�{"&��"u9�E#=1}�}��d�P*�q�26�w�Q��&0X�^$փ�!l/qw'G�l0��PO]���[��D�1��d�����;�B�ϣ v��=�=	r�~�И�6��61m4�-t&5��4�I��e�*8�U��D�6�F��V|<�����R�m<G[y�CA�6��M�2%���`�d���ց��0,8}7�ہW��:x��I3���ΠJ��4ŭ� ��pH��V�����b/�*���`��r�I�B�F���7��ߘ�.�G+�% q �zR0�o|ɿ|�s��~>��fD	�:2׾wZ�[�t�xc��<����1����넼G����J�����ZL�W��/L��[<��s����8���$��N���4#�:�
K��7��iL�N���I�e&?*�`L`����&��Q�H�a��6p�k����d-*F���/29�������n����d�9�a��<�y�K�>�O�T�#{���(���y�ލ�%!$\w�Z��E��=qz���jӍ�M}IM���3��������$/7�o��mE?i5�p��cx���z�{�A����c �&�ԍn��ϩa��'-I���#�v��"�r����&�T!�8���\�z�S]�1���kP8�ך���H��?���M���LC#m�A�4:�vY�^��i�*s�׊#�N,}��OBP���aE���<W�'}����"����B'Ag@%H'5���
Ef"�y���Z�8��>BJ��cf�n6����V \9���L륤�,fEbl�O"��*��GF(/�)n��E�$��o̥�fgfc)�M�RO���H�p�5����~b<�ɏ�s7Cco$ze��i�2�}��xX�M;�r+}��vx7�Z��$ym�迦�l���<�K�H`��W�}v��I�*_2�����o-Q����Z�7��6ŏn�->���0^��J�eF��� �ޢz`�,z�qr��B�@���f;z�2�3��$��L-�3�*m(�%"H\��R�G�C�8�)�� ���
~:rY{�l���ܵ��5�,<q["*riL3F�6&�e\���s1�qE���q�|�o���:tQ�"������{5� N��B��uj��;�M�#"�!.y���֬Ճ�&�9pf��,��0��t�.�-�>�ᦫ����G"&�9�~uWV��7��Q'G�X�dE���$�ml�[��ɚ0�;��ws�Fd���'6�4o)[�m��a�؍t�!�ɖ%��46����_G�^�lgf�A�d���T�kǦ�/_M4i	Ȩ�k�b�V�M ���Q86�	|JpU�-���ʭJ���Ã#���u�ߍ�ΊdYα�j���	��-��Ě�$5�I���zL@��|"�-�:c�E�m�zXN��]�Q#Gm�V2�Ap ��OAB����R���=�+Ѭ���i�V�k���=îF��x�S���پ��������~�?7	���B��M��~�d��܌7�.ƊE�q[DM�ka�)����/;��x����濆 PSB��e�N�W�4i�y+[դ���&�k��vv� �%^y֢�x $m<��~��ڬU��������K��{�����\["1ſ�Ї�1Ep���*�o�mAt�ё�.�K�q�������}9Í7�E]�rW���Xk�V�9����R���$���G"S����v�����Q:�b�E<0��,U�'�\����o$7Ŷ˾��dl%�p����f?/������|R c��W6�N�Û����^B��VP4v���C�i�*�qW����ꋢ��� Qim$q��ח�c�fY�<ЄD׮����Db�rE^u�\p�/6�H�ɔ��l�[�D��Q@�Ez�1�vٮ	����mD�~vk��~2W����'ve��e���e�sH2���2��N<j��8v1Z�=7����s��l+�}��N�ѹ�}O`�֒5�:���|f"�{��NEXP�8��7�cd&�M{s��[
����˟�.!�f4�7Ɗ�ݱ�qgLm�� =��9j $&�j#�6�����#�3K=�rp#T�g ��"K ��p/�[��7��&O���,�:�V'�E"V�A�lf���q�AlDt,���H�dD�D�EU&!Dr;���<�. �r�[�nA��	E��U�C-�+����&Ɖ��@	�d���	�%��@]Qg�b�n]�*��*jw��96���Asnw��}�B9�/srb� &l�mL���i�Qa,%B"�'Yd�>���Ȓ�C2`5���t-v�v]��������W�m���}&j�d�P�[�b��nl~9#R�y�I��P٥�ds"�J�J �`<��S�~뷰���6���^��� ���F��jR
���~w�t�@P"7��L-�P(��V������h\�)0ˉ;A�{��>
�K����� Fe��6d��u�);2HZ��9T��\��d�f�����7�{E<i���9��Ͼõג��,���/�.�hl	��y�d��|���nr�q��kv�������=+�Rjs8�5J�W�0��݌�l� {��^��.�lLM��1�,���[�MFc	��vn�#�"t���G�&��X��q�w/�w~�=Q�F�ҕ�b�Gi�l<���Ɵ���F��lQ�ṇ� �b��A8��LO����߼�#q�=O��C�Jda*��2~?�,��?k��z'?�t����89}�� .p'=�G/��1'�[oK������%�u�F��
�er����9祯�+Q7��궺����ud]>�u%~�	�ݗt��dɒصkWڅ��s��y��S��'�'ѣ�JMX[����@v��bP
�_0'��A�ѻ����‌L:qQ\ĄTf�R�|c8� ]�$�.��u4q�y_�`���.���U�{/!���=&9b��L��Y�~�9A�8&	�\Y;v�E��J}J�&�)�3�[�"���e�1�m#;!���<%=Hk�LL ̃ˎ������kn~{lۃ�}�R���u��M4��;����w�w�0�7)Ǵ��� y�%������>���ٸ� ,9Wk�B̕2��� �/Q�0߆��w��)�\%���N�|oL�s�!@�f���}�`�)���'�%�\�.N�u��:�OBt�̏ɐz�V2c�"A1����y����<��o1���(3ߔ7����]���!:�ג2rc� W��S#a6�T�r �"^��Sc�ԋ�#�}d����a��k��_�Z¥$��!��,yo����"g�n�>8��ɑ��?c�����9Yμb�~͊gui{�c��/`�9�1�Y��Ȃ5�NN�&�5�;��L�)-Q���.�C0c)	ǧuvc��OĜ8r%���Q��n���� ��ς��r1���x�-t���"-��CiFUI�ox�!��ۯ2� ��&{��@#I�=�XQՁ8L.�.!b`"d�UFU�l��{ �)��E0p{������ԟ���h+X
��<`�����8-�`4@�0;h	��r��Y�1�>�J7�x�z��i�9s� ΤLs�J��y�N"R�y5��5�۸�*� �K�_��9V�������o~ë!Ni��j(ت����{s���)	��$�6:7Fo��v��P����*�Q'/����Q��� ��q�|�l����$��V�G' @�Hk8�@�!]���N�r��&�t�>���MR�L�W]uU��2>���Ҁ`��������	lz�,�0��*���~́��$��ƅ��<��S $�Unjs���C�)Q5`)��"ਏ�,#s.W�!���Q,����┧̫�GQ�C��(l�$����� �̪$+�XY�}7��7�Nƙ��GBq��`=��@.܃�X!po1i7�:t��g���4�Z_��h�R'%�Q	|�16F�^�nS*�e1�Lvm���`)T�#KHt:��_��P�?������  @ IDAT�n�	��$'�p�j�L_rp#�ߵ)N���+��ؕ�Q T� \�wj��Yn�@����D������su�G�o5�����HR��]�����)�}ӂ�!`�����[��j���UY�EM��JR����͂��l����G��|�=��x���
 g��lDq��(n�am]L��c�?:v�D�Rn�<�Ց�F�Ύ�N&����7o�����32Ɏ����X>HM�E�r��^�ٹ!�If�
���㔭0:{)\�Ŀ�)��ۈ�1�s�����}��7�O`�p=�R��e]֙��\���kbQϝ�{��~����߆�t�/���4s����pX�&wk��ޟ���h�R��4^�P��[F}�5}�k���cc���c�c��{�F��4���?��dS���.�Y�����wV/��Jx��#���B���d�L�p	$�ˌ���C8�ȷ�"���/�P?z���#�e_?k��ɞ�;�<�.�j��g<�	�&2H�K�A�����^S�W�T�o�pr����=���^��n�vc��(�\�؍�2RH��!-,�u�{@�H�e�@����WfF���^HF�fOd�D��'��c��t�倥I�<��~��e��&b�"oӗ@8�p��޶>V���_\�)��G���j�����3�%�ĈE�G��⎈�ضc7d�;��;([��$�L�l��H,�{IL���I��۰�M8"	W.�������\�͍�w�BV�t�K��A�[e׮������A��L�D�'؋rgb;z�ј�F�u��Ѧ�y�����3�WŦ�vL��+�GY�Y\�\�S�S��UpTp=+��Mނ�"F��+�ٹ�?���\#pU���'���G�d�p'�]�>�B��_�xV�w�#㖻��"���'��,,�s'�糒�Z�F3����6�Y���屬�Z,9ߎ���G?4�!6�sV�<�g�J�>	�tb̰�u(��@�ȷ���A��v��?O��-���<��6	�8��L���}�#�n!�3����Q��Tڥ	�[�}�X�=@NbnDdӋUb-Qqr�Qg0��0u���o]�ǩU�B�]De�bm�U�gGֿ��=����΃��{�c�/;	K�o|C�����wQZ$/���c�=)�n�K���#�1���h�3���L��j�L�1y�tY"!�֨�y�w?랳e�
v�A���c'���yy���'���i|t?K�r�F��$)Y|LW�"�}K��ln]�n�FB�	��Y _+���#����Jcΐ9���5�"�7�Di�I1C�:"�bp�����W��ʽ��Q>-�Z�嬕�
z�z�V �;M��JM�L�@�������l���5�����X���B!<N���&6#r��lxAX��u�9�����/Ɵ����v7��F���y�U��լ[w<���ʂ]{��n�bO"��,g�uV|�����	�r�sݣ�x��o_oz�9W��q"V!�\;F7��U�I���/����4��&N��lC��p�8���
�5)��~�B ���m+���:>i8���:����~t`3pC��b�4ч�	D��������k8u�)
���m]��p�;��a�W	�Ģ���*�V��'s�A��)�Fd�Ua+�\J��9��˵\\�V�q�c��S�/�(��W��U��\�B|=����]��q��@�����d��O�Ĝ�k ��s!��蟼����o���i=D��dƢ�<��}���ƚ�RZD ɉ5%`�aO{sl�їb���<J�*E&��"�v�������m?}��T& ��)ל?Z�	�Ⱦ�c,�aW-�xl�:6��t,�9j�Ԩ��I]�'o������Hէ�*Q1��S�;:���+��V���X�m�c��Q$^{����==�2�(Ee�]�	w�A1��
�O�I lM8�Dm�C1����`��U�RQ��[ańݤ\� U�&w�Lu~�(o�&�!{��4��7��~���v@��=��Df�n8���x�S����;����c�8�R���(�8���BQG�������W�M�0�d���ᚧ�-ę
�&�\O�br�0�8j}�$�<XF!��,�_9�~�x*�/�'Ax����F{/\F/\b��v�����EGQ.q�}K=�T�UPԳ/�g���V\�ZD"l֤	� ����
G:�G��k��l�������8�����M	�U3%D�Z����������}֏�a����q�⼄Dn����\'��|�;�O��Ox�@�a�t�W��#�4XH�'�B�t>K&�� 0zf�����Wr*e��A�c�����;t�c^�n .�pd0R�iω�5OHR������d���0��������6ES�Z�vWl��+1�|/��X �s����_����`���S���5i����L�|���fD��*Ů�j�1�v���梸��[�{W|�UX2�re\�O>���J�)CT-�6��/5~��O����ظ�B���1/WA�a����l��x�{]"Q�끻?�i;���}<O�	w�}]��7=3��u�c�������J�k���_[q�ό�ì�\KP|���eK��y��ݬ�/�:�z�:�0���c����7�T�4T��n�Qa}uz4n��qۭ_g�Х � ͉9d\O}����|fl�
6�e�ncE0����p;��+.�[���|�v5q%r@(�_��Gә*"�Kb��Qt��oȿ�Dw������o����p������O@ʳ�)���H��a�^�+�_�M�t�ɺ�l�{2 2"���:����`}� RE��ug-�p�c(�yȇ#19́J�(��
D)O�yj�0�I��s�bj����%��稧2Q��k��lq�`�����B�����<��ه����X����M����X�(l�+Õ �Zk,��R2B��������~;mP��v���-��s���$�6^�,���R?�K��7��̳"�=D��in��Iw����%ZK����G_��j�~Oُ`~���o�[�p�ы7)i pj���?T�"�y'�J�Qt�L���W��Ա.�`kCP���?�ݝ.���(Yw�y~n�y?$�Q��QXC�̀��7'��`�����/������� ��g��+p�0u�����`�/��4�%�	ʘ�������}�U���>X
U���½�b�O���u�U8�l
�f�;��g��a��U���Em�'3��ܲ���Q�� JjY}�p�۱g74M��\�	����ydf�~��=�<�����k�������4'�i"̎',���=��;Jq>�E~������g~����%�[?�~x��/|abee��$����ޟ�eS���S�/�V��D���
> ]
 �����,_�4ϱC�N`O��x�^��� �,&���m�>�w��DAlS����^��M�)�P%�ܸ�sO��3�)�/�!����UL� &�ڗ
��
ބ������"���8�)�M������㼋��t����-����Bp.�������X�b-��!W�v;���\<WV�O�eW���� �e\�@��G������iq���e���!�e�t$7�=wܷb��2҅$�E�PB���}�=z�([3�o���	t�L��g?���ԧ>5V�Z���=�/<$�۶o��[�%���1>1�?�^�˻cn�h�^�]?���5��������XլX"@��q�߮�3:���Q"�k1B� ���3��~�$��ٛ��}��8��7᰷(�x!b��؀�"�Qko����{6�C�J���di�������r����?����%(�Y;Ew�U��cb(�R�\��(�!�ə����8�x\����n�e���IH��6�YxK#�ĺu��-��e���Dm:�����ʧ"���zvh�%�9��ʾ�� ?��pt�MS�Sr����>U<q]��Gc�m����Nvs*�AR�G@�RwR�	6��J���bt�d ��e���3[�w~�ocb�y���	�CJ�r���`�l=�,V��+P�&N�>�Vt�#�'�M���(>1���禝�2z�J^�-�G"�G��X.Xp�{7!u��6�޽�@|���X���� ��	ԧ�k8'M�Q��#v'��QRpkz��=|f
eUꍏ~�<�ww�LT��7��4s���"F�����W�������n(�ׯ�+��=��
*g�K��2;�6��8_����K�����bz�h�T����2J���('{W��6G/��E87	�,����-�h�c-�׹QiV��b�r�E��$�}߼�*��/϶H�"�J�&Ns��/�I��~���:�*?���-�����I�DW�i�\�%7?��/I�J�ȕݑ����ۈdw�R`B��Z7��)@$*��]�^gf���U�z9�鳒�����p#���ӓ�ӌ
0�x�;R��M��X����N��bd�����ezr�@!�'G/�N�.`T�#Tz�q�~!Z+�\��NkB#��G���wDg˥q�������BLI��4��NbU�H���5�GeN�6�"�5���E�����O��_��ܽ8$��>��p�ʫ����1��ߋ��'�h	bYZa��F����I�� a����\;1��}�\,%Q���P�>*�I}�B�=��T�R�n
	��eP�%�a�����Kb�.��ւ$Pb� �� ?�Ƣo9&R���CT|W� 
����QK��`^%&s����JnԈ
�m5�RC!k��/�h��3�0�18:�ؾ� ��ߗ.]� 951��1m��D{	��cosm����n�
�E<v!pM8W=�{p��֎��u���+b����e�M6#f���6$#BIQ�VE,Qjj���i��Z欦؃�bVEL��YM�<l3�DtΊ����AH�y���.u�L���=�"���k��������M񇄆�W���K\��<̄]�%N�O��Y��l^�������{u�G�O.[�>���Һ�F�����O'�~(T���x����O~�toK�t~br�J�"\�J,��L�
Ĥç���-1t�kb���+��%�kW� v�!A\�!���K��ܥ����������$ZVBO���^Zb҂�cvrzkkl��3��;�F����%�g�Z{v�y,@�wI����1g�qT�'<�����z��]5H+�>�~�� �� $��K���'�g��-�_����J0 `�4�J�����h�_ay�����2�V#x�ҥ��oq��2:>OO�Ǆy�E����y8���o� (5��7D����q,2&""A��#��&��f���09��z0en�Cܳ9t^�HW�rXOMwCS�7i�{b1�c�b���*:H*��l�)��i2.�	��ĺ��\3��|�&G����)(N���D,�5���$�S��(��(&��!SHs��4	�Ip���=qn
3�Yw3MW��^�Q0�y�f�p�,|�s�xOs(�x�9��慿��4ZJ����%�I��>65}Qt��	�����ŏL�}Ѓ}?����W\;v ��!YX�" ^z��W�"&�?�b�p�i�[�u��_O�Na�l��lG���yE�Ȯ��.�Xt��`��2�l�qZ,}�/��ߍ��T<͒�ev\(�qv@�Fc����X�:�k����g<%%"Ƚ���;~������B�QU�i��f�=07�Q�61_�;�UFbՊb�8@_A�����>FN����D,���Z]��H2���z�+㝟�b|�+R���gc�%%�~�{(܉�v$��Aq8�'Y^��N�%s���`�E��+���-��u����t3�}Vb��0�Ζ��.���{��L��{;p�g|o��ݾ�W,�������6�͹�?�	x�e����ɾ5i��� �e�(�wd�ADp���8�<�u��^ǋ+�^�*ja�3����l�EP�aJK��{�6I��%����/_��$.���/|='����ooRY��!2KȔ�! �\�qM�#J�� �i�۰�qT:OL�H*��х�20�|�.��Y7�W��@�ۍ:fwĵ�<XE���WZ��#`�������H�����x�[�ɶB��Bh F�pP�.@�.׬�݇8<��<'T7�� T�v2�3VcZ���0MxB�����%^��L$�j>%�!����cڼ�}r[��F�~����-n�h:��H<Źf�:�k���W0~k�_ڨ+�%#f�ͯ���$�f?����ˮ�w�����3:�J1S�4T�֟\wܶ4<hQ\��b��؈C�P�M�������TK���8�������8�חj�O��`A��o����y6�_��H�={f�N1��ɞ{�w�N$.	��m,�U7�oY|H�mؘj�4��	P�X��"�8�$��}��p����5�j�0�3K�g>�\C�C��,&Z�Rq�� T�s��'����1�hW=��t\��nh�k�~�����*#
b=L<GG'v�������^ud�?~OA4Φ�~���%p�@�^?����Ug�rPWX���q���v�o�zL,* f��y��"Qg#t	I���נTs��n�d���R]�ӍЅ�V��0�~�Ν !;�k3��<�<�xp�U�K�Ԅ"��m5����/�qj���h͵C���K������G��⻭�bL�-����܎om������!��#��7D릙xcj�cuH>���WaC��b:�Lf73C�pn��A��[�n���a�"��`?V���V��!���RD�m����򫸿��n�M ��Y���Da�J��C�}j$��0�*�N닕�%��J���{?�I�,�1c|�h3�lB,�(ˊ�-�a�iF������Z$����<R9X%���z�hK��HR�k�\vttgb"]�Wۈ7"��"9)��G�/�p��?>1=�Bc�b�v/$�<��iS0�5T�*���"��D@AO��9#����U����F_��#E��v�E�y��3��R)T��~�������f��m�ؘҹ�vŊK������N��  ���U5@Qf����5P-��a����}�렵�L����RE �S�{ԑ!=D���G�@2����C�,�WM���&��'���Ѹg�S|0!\��yKHV��#�c���֕?��!�����.�P	�N8�2Γ�Hc�{~y+i�oE�MJ6�Y��oW%1C�	��H����eV�m�a��D
�yƣ��YI.������ U3��,R�W>�l1�Ԍ��""nW�'�ǽpURT��>�EE��IX�5�Jf��~�%�����mI�&��F����?6���~���!�����T�ؙ3�_�P5���_:�+�����-8�����J��.$�HJ�0İ
w�(�nERbj���5�����ϊj�[��z62�e�Ѕ(��j`�F��G�ȶx6�{�.�(�3�ȗ�Q��+-Y�&[�q�2��s��/]�݇�d^sO�D�>�.�0���TIM|��9�_ÅL���9w]z�
��������!}B�:m���A��ź5�&��?c��p/���
0i�O[+�$�L��	{�I:��GuT,X��yW�._.�9�S�c�Xҁ���j���#�����?���[���V�ƸV_;@����sW�t�	�onݑҊx��kc&jE5��qL� ��9�d�U:��b�4@����h���B �u~�L"xj>A+�ϓ��Mz�����D�B2���s��b��[��h�B?Ϡ��D�"wVA���%�_����?�
�H�̭C]{�+�����Z���Ϗ��_���a���R�.����}R��L��+Y��O����i2j������Y�t����ׯ�=7S����U�|$&eS�7b�%Y�s:3>t��x|�3 ����# ̵ ��x�-l��s8w'KcH����d-���x�8�N̹��R�V¥w�{?�->��T�CU��x�DQ]&ފs#xs�o����=�疳�����t������Sl�L��x���P��@���̜��H�"�[^?+V>�w���jơ}�+�0H^{�G������ 7t��Bu�x��P�x��÷ǒψw�����,xl(���pȳ&mJL	�X	E��Q��s��!�r�<`ȣ��_I=H��Q?9��������I/Hm��*��6,��C��.�r\qſœ�O�*�����S��8��fC�D��!p��D�
�^|���h�����#�S�2�U�����DL��n�G}4��� T4o�_T���H����0�?�@�Ey���ف�j����݁�"C5.v=�謇  >+��^�$P"BVX��2D��� ���7��8E�"}=���m$]ϧ�$����D�"1�����'K1��}�~�Q��1���Pek�X�^�]ì�)����/o;��w��^��[�-�%N�D`�ທ�߿�=�kY���>�D��7�����ݰ"���߽����?Fz�$��rw�q���\|���­I[H� ��P���� ��v���cִ�x�Z!j��h�0و�)	IV}Dcy�nPs�E=�b�V������d"f�vww�C=!��5�>	L�QwJG��V��?�eFT��4�?�U�Bi�z6-+�\�OG&��`?�X�Z&�g�*�dM��x|y�ob͐`� �w�#'�P
3�)����{��m�H�S��Z���峐�Vah�Ud��! T1":k0�Ύ��Y9w�v{ǝ�0����&�c�^��3Y���0!�ڷD[���^*�ɣ�5��p�Cڠ?Hu�*��P3ɂ9Mq��fs��8)�j�5��u=����F�~?��J"������m��R��{����	�!*�'�����9�w�����(��3�M��ŋ�u�{]�X%zc["&�0��߾����K��@�N�i���p��o}7f~���{-&��v�d�0z�S����;�+���a�1i>��L8�ө�����L�=e�D��Rg��#1����o1آ�w�"�p����4~JT| ����ZHJ,>s�D]��� �&8��+M}l��|X�m95�9�L�5㊭�e邒1f�m����(�*އ����Ƣ���@`_g�ʮ��D)b��ftM�|� ��� �I�;�P�';'j{��|bV,�Lt+�L&XF����}�)����b����Fl��q�i'ǹg��6Ȯ`��F� Ի�bӈ�_�z��������k�-�f���V���?���3��˗'�KH��ҵ�Y�fe �v,�x��؈M�q#R�v�>$Iգ����_�N�� ��Bw�� v\�=���G,>%�!�+���k(;�Z��c�8��{U�턃�7=���ĈE�3DV.v��r�ʡTXC
e�����#����~�S�@#�fz��Qc�7�I���M�$���n�m���w�}䗜�d+J~���,���T�?��?��{���Q&�ƶĴF�
 �-q1p�#��9$�EZ�,jqT���oLB�ѱ��g�������v���??1����;�/���髄�T\�ͩ^I*{�o�\#~�������^���Ko�����H��
�6��_n��~eI���W Fŧ-�pl@|E�e	"��nP�W�A'��O�:���'�h��v⚔��+$v�����M��A�rXO<{�U1����A0��F����9b��%[D�߾��L�8���UX�x�����tC������֭��>-�m) ��HF*9�����e4�ʙ쭹3�S�Apx��=��A�T� -¦{���8�ԂD�M��d��P
����&�nR멆�T�s�W/Du܎=�b��>.��D�Z�J;R5�l����Y1������a�X�G�!�P� ԋ�WUi��y�[������l�������? ��p;��R����[��mKl�M�JQ�9h1� �sQ�ׄUd�KT�
Yן����G�v�Mhc\"fq��CE*���E%����C�2E5�F�3^�j��Vtt�3�뛍!1�w9FR� R�����V��|����2�Ȉ=چgrN3̄��i���\'	f����I�5Q�Y�}�߁��`���	�iؑ1�M�]/�G?��4�ε�J�&ƕD����>}O&���wG�O}����-J����?��v���$_C�flD�B2R:N�B�!��`v�Z����ЀM����|���K.N�2ގ��xBb�J�|�ҥq�!��8P5��TCD�Ʈm�Sψ_,�. �m�0���D(
�IeDz�����&�<Mψ�D�Ł�0����q��Q�v0a��6 �{���x��<��RD��p'��rv8p��IJ�ͼLy�M�:���� U�rV�t��8���3�$�`_5 �0G�{ڔs���.���,���+�0D�G��υm���fE�@��X�A5�u�uncASuz&���٪�S�t�x�*�QC�HG� T���s�Q3��Tm�{&y=�����R���i��Z)�~>("d��!l?����e�AA}j����_����[c�Vvm����f�=�J6��� ���Wv_�8��Rs����x���̷���OG�rQ���8��J�0�V�?p�E��9�kQ�haݬpW�=_U d���-lKF�Y���OX �nC�u�n%�F� ˄��!��!��uG-���H)��1�>2��H�C�v���JOJ�b�!���*'n�\�M�;*EX��8�l���؀H��9;$�����㱒�8����Ӏr�`,,��'���"�^h�A��0�"E�k��2n�ց
L���v\�-sr�&+���ĭob�<%(������MB�T�i�8�o�9�S��D�g�6!1a�Lc��ڙ�8;~p���?^�m^�	��x�P����~�vj�=��Y&U )��&���vLd�:��[�~dJDtS��-\M�
�M�2�,q�m]�0�����k$u��GUDL=�+�� 
n�U�Z�:<bS�0Z;O��oX�����k��m��M�Hd�Z�Xm9�§��OR��O�U��H2#dζ�_���*���l#E)��X��A�9��
`X>���:D䖐&j�(��|5��u�G1a_�6�EW��۟Y)��V1WUq�z�{ֲ�Ѫ�f�Nh�)����iBꡐ2�/�5�B���;���⨎J��=�X�D4�͙3�ER (���5�`��B�Z_P���H���dS�gc���h�<�*ǞB�s�9(�r�dX�T��-���,��2��^�漁���V�tSF��o�,�Ŏ�(ZQ����A��P&���(m�rS8ģ��~���� ё��c;�$�q^fgo*�Ӱ*���H�b?�I����Oa��x�z�q���0�9=B�ꈆά� �x"R4H��� ��;CX��y���)Z��1�ed�ٻ���_�~ȼ3�@E��H%F?U�0�����A$|B6�뙸4�L��5t5�׽�� <�zک陾KxP��&$&^,$�g>�%�m}ҕogOoA��}��`1^����ޟ/%�e���۟Čj����:� 6��(~)��_�C��D~8���b!��͆�q��-�P݉d�NMѯ�}l�z�P)ՙ�
����:�����;I+A�J�LrD�~��p�C�u�7���-�O/�߄�Ww����J���=�<5�	K`��bd��I pN�F[(�#�ܦ'�k�ob����}�^"� C��ZM{�]؁���f���_��S��0,Ϟ3?��51�o9��� Wq+�hGt��-k�.������,$�@����[�EC|�ɂ,!�lF�P�SC� )b���m�@��ؒ�MqJ
Hu�)'�m���|ǹ��t��]��[�3�,,2)}3H)D�!f�n@���\��B";�"�ӄ�W�H)�&���,�e16�����bO��HVm@e�,Y�M��6�j�1I�&�\��qGSi�kv��X��)AQ$s���Cİl����z=�=9����B	�yT̄�ȱ�I�
S��ׂ��W=�?�0{`�G���-s[���@���wc�$tJ�[���f$�{��w%"���SwRb"��s�2�z-زdɒ$�Μ9�Q0�yV{�i���}$����I�[Jyp���+U��0/� �
���:B����D?kTt��G���ݗ�I!g�̦vn�=�G�?��j�G�`+H;� v=�B�oi���~u�jWK0X\H9@3���������xW<���\��3��y���`��8~�'�蠎�I`�ހ^v6�&㵩sA�^APԾ�#>�:��
��C�����Hݬ�GӺ��.�B�	� � �H?������X��n$�[3�Y��Da�g#�1��E�Fd-�5�>�E�	��-@��7����X��Ul(�\K�.^���up���o�	�����mmnт{���/��3:��a>��FjŁ]]�"^�?���/M�Ğ�#YUV e��8P�p��0܊��<�k6<5������zb��V�o#�{�:������!&F���8*V�Y�����_Q[N�%�E��o��i�L��3A�y�fޛg�H[�����z% y�MuGºA؉l>��X����y���e�d^�?������O{�M��$%�FbL���]�r��'�t��2U+|�6��HP|��G�^�r��d�7����}D�����]���s���t2�-�{�w� z"F�sX����S��	bр˲#c^�A2��v쉶�ӱ���Ҫ[��ѥ�٣�9n�8�y��UR�~�n��}��B  �~�����7L'Ŵ=_'��9���vG	c�0�%��)�)	�"�zi?z� �C�1�����Z��_?�:fơ��:��m/J�ᘣ倨j90j�A�XK�\_����eE59-�y�L�3]��{H�}0����Һ���?�����#f�������?x n���+\�d	���;|�!+�1�*b�2L_k�R����6Qo���A\�uq�O��X�׺'�u�ݸR+�{GA!T�j%���V���{�|q,h�C疑D� E��i��6���ͨo��v$�"���x��#j��0�E��I'���l���D�㍨�
R*��E�^��N�Wɬ��N�"jã����m��I�nJ7Id���\W�4
�����o����q���1~��gyG�
iX	�g$c7p"aI�Ef\�G�� 0�{��
ፏ���K�"��W�+N�������M��2OC�����*��s�d"���7�`�2o�%�R���-�7ӡ^6@�I}�D8c����������8��?A��U�l�-�X7b$》��fw�>nB �A$��#XE�:��{ �V����)UP�1M���@�k{�7� ڍ��1�`y.��1c���H��O~~I�v��h�Gri��Z$��3e4'}x'1q:���U ��m�e
A�`��T�n�p~g̟k�$q3�h�t���v-���5��{+D�IAd�G�|"�|K��98��# ��!̑9OnB��y0�H�{	>b��^��hb��w.�$���0�bLo%����N3��(^�=��K�cl��Ƭ�����D2�!� ��6�?�ۗ]?��[��z\훣{�jT.�7t��g)6�����+�0�zrs�Q8ڌޔ�ͺ��.��|lI��K:c4�޿a60{ꙧc-��T 2U�*˸�F@��_W�X�h}��c֐�j�r|�!
G!���B5a�)�����Pe��~�ԛ`Jc���H��������Ͽ��KƼǎU�+(�]������.�,N:�4�<T{�TmRb2�&-ƾXK�׿���x����AL�p!�'���& �s�_��wNl^}�n��V���f�o�YB�Fl9!������Ku�|\�#�$S�@B �Ӏ��w.�YdV�ܡH8��DմC���(.��i٭��>�wi��p��(�z�vԊ1p(�IcE"�~�I�=��@��L��랖���2A$|���Jo �ۍ��VO�'�Q'�O�s�LI�8��q_Z�&����@J��Cc(������8��cS���zTT9+]MѦڍ��� �ST]�	�Jt�M�K�G�2�ØQGv���ǹ����]M\	ۯB�J�J��ԑ�����z��k��H�4�k+x�L�( �T��
�uK�ZU�4'JU��ЭM��N3g}�>m�&�0FV#��.���Q��|&�bon��A�8�!�g�VP)fG�6����0_ym�ueF�]�³�q�FQ	������~0N?���/fd�ML$$v��}�K�w���d+bȡ�F���ސf�yt�����8�bbvϖ'�o�}�w	���0�1�t���<K�] rp�N+�P�j�	S�GJ������4��m��ħ��߸�J��D�b��>�k/Ȧ|"��������B�H6�3M�o� 1�d�M�M FsatE����WBh/�h0��'�±y�+��#1I��=JX6��=��*�@�Hssj���S����A������_��.���~�D��b8�����5��q��r���?�3:��lۀ�
/��j���%�c��=���Y?��AK>k!bދشJęde0rr���<����8Ӕfq��dLF��v�:iSݓ����Ϳ>���=�L�\,�u�6��Lu����6?a7�a���5mS�Ο�w,[�,G���n�w��H@�b��� q����7�������SDjr#�b�%E�=�:��P�}�b;a����gb���I2�t�%�*,Uw�/A+:&�����qo-�n���f^4P�kŚb<��'>�ornm*���]��C��s3c��*������G�k.�&�h5�`���AU3�U���"��|>+=��S)!��_�w%��y��=z�gB?�A�DC��3+��u ��"�"�-#�k�k@V�qi���Xhڜ��o?��8��R.���l���MQص6��7��&���5qǭK���yd7�-���3B@�`�Q�ʞ��ؘC��h��!rr�j�D'�OiJVgĚ${�1ǧz����|d�*�ǉz���H||����%5�8���w��biMǾe�}S�l���{����ɮ��9C��{#@���I���moM��ӫ$��3b�H����t����^��߼'��δ7q�z�C��-d̺��E|7���R�Wc�8����㏧�YC�����^�P��pO_C-J�s�"�)L�ل��1`6��ۃ���_?���=�_ �n��V#-�t�� B��-f���^�L����F� 2�FP��w�s��_��H�I����O��Z�iMS.������.E˂"C�E2c����AR-}ME�Q���0f��c�&ţ���AY�B��0^�y�!p5���*P{��YI�c�A�	�$0��ʹ�����"u�'k֝� X��T�W!^�C0F�zu*�Hg�_�O�'���:Y�ʦJWC�k:���kn�K%D���T�H�"1`���HX!�I����4ɭ���EQJ��y�N �C;�D-��	�N�b�.׍!f��&I��'x�K���?_"1�)��-�m?,Xn�n-׬^��S�F���b�nK&�{h��}���W_}5�_�d9�`�O�B/�0����R�a/��i��;;����5mq�Lg����Ӹ^��z���}�i[x�.�QIC@��Q���wd�����'�-��_D�сx�y�k�&�(!��f`���;���?�����Q�:��7m(6G�Z� �kG��:�?2w�wT��T��
0I�I=�c���Y^=UsΦjmY_�9�+����]��6V�HC�7ϋ�����s�FW4�  +IDAT/��t>;5�;�7������=��:�/���Ϛ�)/�LZ��y��!��M��1]�`�o��]�~_�pa�|��I�w���i/���{��N5��k�	�>j)�t��tu���)��[���5����|����%�{��}��+�����1�d*��'�&c[��cx�~�E�x��1�֮H>~��f<n�#^g~�����G0 ��6�Yb�w��?_̴����K!��v��X�(�L=۹$Bs>��Jb4�D��8a�[N���#��n��]�}���xv��dE%��m��������uF�Ϸ+1��(y���8f��u�]G�j*i���׽XIzȘ^6b�3%v(���ڽn&��2�y;_�T�k_h0>7�4''���>q�_�D�m�f`W���������{�� ��#�����������C���O|��9I�Cd��]2ď���}���^6b2�Dz�����㏧����:+��A8X���)⻃�~]W���M9!�����M�v�_��s���Y�V�JM���SS����}��xxOL��WdK��}�o�2V�t�~	���� ;��
y^��-gڎ7������2/1ٝ�+I�D���O���\r�%�f��k���!a�ڜb�γ'�&˧������{
��b�"���U�x�+��xb�;R����<3��֡�a!�����Zz�px��&��H+x���JL��L�(u�`䒉�I<�.��Ҥ�y}NE_��_� �RG�����kj9/��=�w;�ɟ>>�f<1y9���o�ΈC�{��\��J�V�6���G�����G�    IEND�B`�PK   ��W�6U�o � /   images/b829761f-344b-4f5b-9b94-abe91c4d6d49.pngd�PA�.� ������	��?x����������%�����ɽU��[��=����#=�U��(�����,#-���O���y΢C��	P����"8��(�k�X((@����@@A�A@�������/��?t���̓��ZH�<�����yD��m��媥 �k�h�hl�hb��i��_T����D{sWcbO{; �� �!x���)f"%�/��� ���2����91'#3#3� "111��������4��	�Z��:�21yxx0z�1:�X2����01�2��2�C0 �\�= d�M�<�� Sk'WkG����&�n���������Z[�?K��q럃L��abadf������O)�����?���d�g����o_��?��oO���UAD~��;l���;��2�"j��gRn�/��o���u#P��9�8��G#p���ڼ����ϡ�h�|ca�=Í�ai2�B7O3�a
#M�v����x��:~w_|�}t�/�0�=[.V��5��m/s/�oWy��x_����UWw��X��������M/�ׇB(�k-�#5�s-�����Ч��7ƍ��2ط�X��6n���A�M�31���T������c��a
�����v�9��7�R��դ�b�7�h��/t=g�Tg`|ԡ)��ѯ�:�v3�4������?|���7�֏ b���S��K���s��'K�B�[�x(�Љ����{&J��7�4��@�����MH֤gd������XZ^֜�������f����@U��$U�8��+��E�� ����:�و��fi���e>V�x�=E�B#�.�!5Bp�45R��s� $��5��o"��0j���%�%�P��<K_DF�꿅Aj��L��~)'���e�Y�A*�IVL�f`()����q|��,Һ�¹�C��\�,HZ^%������N��/�����AmY���yこ���,�Q�f|CG[A]Y�J�Ӫ��n����T4U-�q-���� ����O����=&�Nd�f�Xq�v C홗cAQk�c�)F�}�o��E��7�>��G��ۭ��A�Z���F`��DÛG��l�j�� ��?n���L�i	݃E�*�F���#�y�K�ys�C�)�l��}��.�� �;��~yYRj����b֫��:���\�2��DK�:Bs@Jo�vp`@�M=���r9�60*��x(�*ۘ$�SR����ȋ1i��&T����B]���Z&}?��͔�?�v�t1"eZA'lG�άI˓��d�.~b�'����2�v�֛�t*�kjʒ�I_5���@Qо0��r�͇��!�Z��ó�[+{'k:b���v�[�NG8 p��J���r	tW�$O�q݅�>Ofp��$g���߷Ο�4+�f�5��m_(�,YU68h�L�F�����M0Ɲ�[�z~pb����|�|�X5x�Sg��ی����&[�02)�*Z��r���S�FO�?�����`)�:����쾣�B�:���8Y1�4�E!���<��������v�z�|іC�f���K��85{�Bz������{�m�t$��N\����mn*�Ѳ6$��[eGkN�"��6�D���~?F��\By[���y��Da���&��5I�� Rs5�G�\�rQ��b?�k��B��͞��Wc�M���c�]�@9��:Z��]����	�\[�?��Տ	�e[T���Ⰲ��蜖Kph��W4�fm*�f Vɸ� u$���k��.^.k��G�G��ct<�תP �͈I0~����`z��B��~��Gj�3p73S�N�:���+�K`�"w)NZ<��$��e�`�1�f�A����J��� f���6^i�QfR4�XXw&��g�`$)Q�Ï��Ƌȼ�Q���dh@�����'�ȝ/"gX'�| �CE�m��́P߯\������c��{�燚�[��Zψ`����Gs�S�k��~�|�xn���A��2�aP��I;����A�ȇ$j2ǐ.�
�9���X����i<��������qQ�N#��zo�Q�V��ws��%̝.�[�}J�դ��x���I�[by�Ĩ�9FM�J~|Ϲ+�i�]*�e��[�Ĩ&$.� "�]燍��X��[��iQt�\�������U�϶�ҰF��Ա�]��Teη9g�ë�����T���Na�۞_A�Ǟ�2S�.�ӱ�r���`Tj�B�j�@Kal�أ�9�4��-X>[�(u�����t T�����1�o��?Y]���S�-�A 8x����aJ�������1,,���9*뀤X�#y}���նP��MCQQgSSmY[UUWiA��j�+����J��3�ە5U=]�Ptje�����×E�i�-�<�zu��Z�������U�b0A$U��gP@S�^�1w+�`�"#ȥ�"4�jkK���^^�����0����!�zd������`*	{�� "�'��������R��n}�)m��#����r��f�様�� �hê��PN�2��U��m5j�����rY�*���gsm3�=y�}0t-Kɐ��/��N���ݸ�w66&UL�-���DY-՟�f����+�ڌȮ�i����)%��?U��%���..B�5o����G�3���JSW��Mr�7y';;x����X��둊\]��!-�S[���Lw�-o�jO���*O��=����vY��J��(�q2�V�B�Y�<zw���� %�v2Z���#15�8J�:�d|�.���s�����JlLö��ƻ?�:��Y������i��t~o��C�r��w"��n���2y�>	�- ��P����~�e�^*)���rVMi�����nPY�UxjPIq����� �����Q))X�MX�&ğ����n��@UU\LfA����E�������/�LJ�U J�I���~��-A>���N7��=rm{�S�ܣlC�󱃃�����ѕ���𒌛
<�z�a�3��?;;a�����,I)x�7�vwB�m�B�������8�M����E����EWi)��ʊ�*��ͨ���` e�H��s����:Gc4Ya"}�hp8��y/WWW���bK��U.��#��G;dg5�P�?<zz��7��ԙ�leX{WgG`it2		� dddOg##W�W��	YC�t66$6�$���P^͓������q:KK�*��.ޏ����J[a�ў�����t|��
BB��W����ie�����~���+������o:�v�uNz�%!2��l�]�J�R����Swr��ʯ��˷3v�pp�Ȅ���d�����[�i6 ��LE���b��1
p��/-��@��UeY99?���2J��s�L�!�88��b�"�Ӕ��#�[�\{-ݴե,�g��:B{�q���*�H������%t+��X�a�KeUx99XY���ӵ�R
h:9v��2��vz���$P>�'-�j��bb�Ź�o����T��N^�	p�4X}f��c�HB�@oo5O3����s����"& ��[��<hr\�������y���@�ep1@.��)�%\
���B�<C�
����5�vG��e&_1��h]�85���]��!�j��g�b��||b�n{;���v�8+��1&&��Ȣ@���;v\+8���T�c{�+}8�O%*	z�#se	 ���td�~#<�VΉ�[QLx{��h%u���ܺq�[T�����9�Oc�]�ۿPdi��::<.7kkk���܃5�+�pJJJ�+UU%�S�;�	G?�s��C�8w;;��|�>��������s��T�(��v�Tɉ[��m�w��{7�,��%����_Ƕ��%Y�j��h���i��������οñ���MM��jjX�eBvW䏡e�6M++ׁ���@/��JG+h�k�7 �n�Q̅֒B�	p�H������y
������8�i���`w�U7���V����]�=�]�����.e��

"� ��/�J���Ve={S�|�aCK�;ll��v��>NʫtJm�Np~nu�/��f�xGui��^��k��M�_��yW 9���\��Y,�SKg!a�caQ8�����o��7��yX89XP3<�j��rT��eYӠ�íf-�V29�"Gs�����=��DN�����kU~o�/j�����LV��k!�i 2yvv-esj���/)	����6��=w�_�*w$N��9g���,~��Ʀ�
�B3_���|p�Gj"҈9�<\:��Bp|Ie͸2�}��������6(���}�%������� p&����7� B�<ul�4�p/m���pNF+]$�ϝ��)uO7S�l�m=I	E�[�y��&�&?����i�}�@�41��}��Pgɳ=]��R�� �uTt`V{6�syn��/���C�G�ߊ��5�;1ҫ�O3��[X8��ԪZJ),8�0��d�U瑺_����R;��}| /Z���&�'�� C`��|"G������Vzl�l��v�ܘ]��l�J����H����x��4-`����Z���+:2ѳ�����WC+����1�w����������O�K�K���<	��_�ρ��B�޺'R:̷*��!�񣁽~��g}3�a-�|E��o��3~x|�FNG�:Fp'�\]0r��b�w�W¦b�C � �ե&-�e�0�Q8i�7ֵ5.R,�t�y���a�W&��x����911t��d���ų�'��������黿�*̐�n
��C����iT����K�̮z���>�kU�6����[�ڄ6g���>�|[�{���0�����ݦ�T�Jz�!%nz��V���^��v��)�ozXU'u7< ��9�q~�Iٟ�5on�e���ы^��H�����HT��M���G)��<����Cg�M��`n92VV��-�{s��hi�j�g,�u��H��#�r?ӿuq������c�ߣ��+f���Z��PF����B!y��pQ�﹥1���%w���Z�p�L�1�|~���?|7΅�f�c?^�_��L�R�cM�4	�9�������0���j�bFk�� $^�]�/[�ᧁ;�G!��	��؏^"���%�L�4��"^Z�j�6�Zf~��@����"��Ǭh�q�f�ҥ��X��g����1����M��R���Q��À��7��*��7���X}���)$� ?����2���WC���?��u���{'�sO��ܐ������ �T��E�+BM�7Z�6Lu���z��Z-*�R�(�%6wD��\��9b���Z	�nI�k�/v������	�P�(�Q�m�JO�����u��T9���E��A�����)v�fQi~��Z��;t�0�!���4�o.Ǖ�ad�p{<3H̛�O]�ͪ����K%�n�m��o��?\h���E�.�Q��a���A"�X�D��G$��;�qcUl���㣫7?�&��I���<5�ѰwQ !�b��з�_?���|�L��*(�Z	�L+2i�	�LM�/ 4�)�84S�RLV��-W������d�����]�#M���ܞ�O�+�ŸX9�e^7��� 9��e�R �-���� !��m�	a>ߧ��NM��3���!�G����'���CϴB��c�#>	�TZ�RiX6ӕ"&�&3戭JY}�$�*�jG������t�s��{	ȢTiG��(M��mn�<�wsG_dx�C{S���6/�YU^�#���{�"��~��V�Ѩ#�0uq1)�ǎI~��MZfh.��%���n��\k{��$p?��N��t$\QB�8oN��׮B�SCw\�v�si�4���M%����	��/c�Y��~.߻���Xm����G����AF���y��'x���9�D,�E��P�iVN��i��-s+-�"=�ϭ~��:�2�����t�}ӯ�H<X�Bc���<�ښL��kσ��5�m�v��Y��OT�՗Y&�ŝ����A�'�M���7x�0�f��e&�L*1"�~,JD�>n�9�^��/�TL�nw�L�,="3�ك<zX_K� 4H��e�^
�@�:�юn�k:��:�9<��M9�]�����<i����5I�N�"UiM��ɉ�ӓS���X�c�k����tt컘����׬잕i����������R�����?��N�G`��h�X��5J<�D/=m���|�u�j��3���_UE�n�B�T�^5I3�NV�W���Tᰢ�]�}����4�A�����2���W9�T�	���+���M s��ێ� tri��de1������}I2 Yg���~<�J�����B����N����F���<�B�\> 7�c��+�CaQ��%�}b��jV�����xD����r3O���eY�cN�.��	}E���zgH�-�#�A}ܨ��]R�2G�.���/7w�o(kC6�Z�)?k���������쬳����lO(K�o^j�Ԉ�+?��f�3���M^�F�a��A=F������lN���4H�������br�z�Xs�%�"����쯭�MB'Z��;�TY�Dl��ݬ��l��e֜��
�O�Ю��f�T�؇Y�,�����܆ĭA��.8�%n3'7�s���W_�ˀFi�����x�%F̰=.��;IL��~[�Z�	������մ��:fķ�ρdj�}�U-�e -)R鯘��ٳq-��\���*٧|���*�\���JIJRl7�I�<��}E�!PC������mjr��4����2��'\���m��z)�p1��g�Q��-�qU��,���
r���4X��[�̱)GK}ZbwԖ<���6W��ϟ�q��|��n7
�{^��:�]�$V��eN��]܉c��#�ji ��1��uB�y�[��`�GOצTw��e�V������7ʿ�לJ�t�5����1322�vX�9��~��HI��g���B��>њ����:��@��ab5���n����%b\"�;c��)i�a�z]IEy�(RZv�G�GɢO��r�q�����^S��X��ӦW�ZI6P�7ypL=����1	���
��[�������	�9�H����]v�L�N��J��4��J@-0�����4y�DY�˗b�Y`����ΊgQy�Rp��O���.������Ña0��@�'���q�9M�M�<�C7D�/ڇ:<�Ԃ�[�+�j /� <C����*���|]�;n=�,���s ��W���������\,���4�l�(�rї�4e�k�oލ�D��ů���_C��wpn}���r�{I�u5yձ�X�c��T���)t������p�V9�c��+.��� �%.�����#�4��0AR�Z/K���9]�, �]F�W[Tk�L���p�D.���J��kH�d�r6����0�þB�����n��y��_-�Z9Ժڈv��d�"��;n5�_��"�2��<�iS�@�d�J:�uD���8��
S�U�5+��;��4���g���HyTa�(�fl\�����Ko(��]�{��&���"c�R*��P.��4P#!ͧ���/�i�o�5;�@hs���5����9&���IYY)ʀ�+w{�9N��z.��ܧ{n[��9<�CW�����*&��8d��J*�v3�9zZ$`�0��93@�̥c|/% ����[p�(p9u�K��o�m�J19�V�����*���5X'�9�$ x�Ԙ��=�S������M����a��Y����py̹��z��\R�Xz�O��0$˛4��}ڨ�/��4�e-���k#�Sț:@���Q~�9�=��������F�?R�`��J�{��t�5��b��%��(�$
*ԙ�6w��&�\�5���uDH?��g�2 햗�lcdA��
Q��ě�%�\~A�`s\�D����	�q��6!_j5Q���]ʚ��$��[u?��bU�}���t�� �����խ��X7����:��h��d#,��Uan��o�.ǖ��q�v���EuTO����oO�,�;�Z)��Y&by�=g��L}8~/����J�$�'�'`��%���B�F��5�f������ �;q/��2��:�gN��#ª~%]2 v��X4�
�����qrQ1���4�'a$8��6IS��)QEI�dq�%P�[����ON!j�������h�؉�����	QD�Ћҽ}��/2�H�"nE7��`�m'M��6�����xg�`�Q�V
�N�nCK܇l4^LyO)�m3<\|�S$P��K���}��+��1\����|�D���[]7i�)�>0|*}��K"t����=�����$C�v�_F���k�8�����{>���iN^W���N+W3ʪ�4
6h_�߽?^.�H5�����w����׬Xd�X}��8�*��W�r?�0E4�go(�f�h� 7�T�7-�-�����$�V�Jeˣc��xg�����Q�M��������(�eL����<?z;zPZQ�����A�);��-2咢N����sK�QK~��Wkןn��N:NObxb�Ѩ=Vj�&�SG#�R���#Ea0��m�{�@��u�D���*s-���v|��h�_�@F��0���[!����?�5&����b�-��\ؒ�
�I���Υ
H�!h��������S��\����l����3z���y+�F,Vȯi����ww�$�mۀ��Y
���il8����K��8&72���I%�3;�
��Xrq�N^6^��<�-�WH���]e���U�RI�������[ǟ�2��-mbT����(Y�nz�C�/	:�eNΔ�TGE�p�l^����ǧW��Wm�F���?p�1�fvv�Y=�+mC��-��*�AӞ*J�P17�l\8�o��B=ryI'��4c��O�Ni[D��dv�U�qy,��F2S��+��ʝ	HoVI}Q���]}�蹞�ŔT��=i5����L�P{�H�"�\���x��������x�h)G![9)J���UaG^GO��"=*�?jA+P%8j4�3�zxD�[��эy)*6u߿�*���d���r��	��Ғ���.-2�kZ<Lcތi~�10�����ݔ����2���z.c�˖�dE�P���7F�����l��[v��	�m{�������i�6��7s��tjѴb
�x��%x��wS�r��.���T�3:��KlK5��q�LUX��ĜH�����o�w	�p��6�Re�l����@pQ9��N%!b�,,��I�z��6��M>\>YUVېJ�_N,����<�x��ڤ��1�n���@����w��|#i�v�[p�'��5IW|d�5�]���g���X樢�R%���6l��DnP0X礸QF�㸾�ge�;Uy��4�NDm��@VnL�f�s����ΦQ'��:ȶ�D����!4�V�(���)�a!��}�Q�*�DW=Ih�_�X�����
!�RK�|n=��=����s�������w�.�"M�4E���B����FX抶F`���9'ɐ���t�wv9�-L.:�w�#�F-��]o�ԅ�/�U��6S~�t)$Y����M�%�O��R���'ڤH0�ι��%?���x8�v �r`~��Tʴ�S�t��|�(��*bk=O��D���i/��ċٟ}�-?���T��]�|�q���Nx/g�E`{�w��W�w���q,�'˶�du�V��Ǚ�~5���E;B�����/$�1��<�.Q_��o�e�,�a��&���4�'��
F锟B$"q�6��0)L�-�v���U�ڵ���!�&�j��ps��k:fj���۱��m3�j�5�Ѫ�'T�K�PJ���O�q������hn)2�=Z�#F�5x������r�9	���kuGP��,_Q�5D��a���*4ʃ�Jk��Ѝӆ��f�e�3>�VhZ�Y7��WB��X��~+=H��<�6٫���r�lx��>���=��`a�da�vuww胰��{aZX?�l+����_4fuOt��EM�����iKS�>4a�ihX~ub� �y&.��5��O��N�A�ͧsB����d�]�	�Yt����@����L�m�X)C�B�D����W�b5�=�_o�*�2�s�wYX;��f��D9b�\ �c��Ě̌R/�u�	�U���M<]�9�1��N�o�X�MIXR[� �����d�qԎ$�r\���D�2�p��a%�?Q{�Q��`�c����W" M0����K �4:�J���m�>��>2G�߫/�)MKљ���������.�ꙭ֐e�)n�쌠:��$t��:Gj�hDs�j,�Y&��(��Ɔ��7gl��"��q��!b��U*�������� J�l^k|
�Ʀ��J�H��J���#�nt7��
jO�*[���S�YB��N�����4�,����u��x��CA	}ٶq�Hxh�$J���v������@�r`�Ê����]W�H�>z����*�����$�s>��C�P�/y�ɞ�Vєp.N�����!��]�������t��+gn�Y"I1=�����7���v洑`����5B{���z�Ѓ���3��=w��fr߸��z�_����|���o����/!�$2Nb��d������?����30|b���?�
cY�2<5A�����3�a9m$��A�6\�5尘Ml�(/��x��֮C��wV�� �sPyu�YFp��w���Q����p~��f7[����~�c��{�jWG:�����������r������(J:�i���>�%D�~2�vN�4��Ë`�S5�����つ� �(���Lp��K	%�A竓\���M����w[c�iQ59[�ӳ8�6�c߼V��@��hn8[��;'���/5� Ļ����':�b��y��_�im0�a��㫳���3Z[N'{�|ͳañ����f�k����m�%g�&*Hk$�����|�c��v�m��fk����Be-uƀ���4��8S������]�r�� C�����ɨ?�$�r;++�3��,~����3������Û�[��W(�u"&�YZ����G�*�*�Z[ŷ8����R$��gjhZ�C��RDБ���6��t8�����H�
��'Ad[�q;�zn���%������*�6T6UZa��������� �*eNZ�8�o�,���9ׯ��c��$2�v�����6��m�~�f�q�K���F����v���3��J�17_V�������v@dd���J�-�r��:�W���O���6�������m�6 �E����P�3rZ"�Q7���3���y���d��<�2Y71�@�����T3 ��B�ܳ�c�.�k�Y��]N�j|_�FKk/��Y�5;L^���Zp��L�j"����f���@��n2kvW�8!��2����͓�Az.�q�M�57�*8y\�غ���iݐ��2)������mgT����%g�j$gp:L[��ھ�����,��6�j{��=(����YK�-���|�2�qX͕�B�)Sr�����2ٖ��u�n��_I��]ܡ�^G7Ӯ���K��"�<TA�̑E^L�U6{��/xȗ���l�o���y�m��3\4�0m��t~͔�3C�a�TE	����ڙ����C��gL�/���(��T���q���qo$f����ͱ6�{=�޴-w�a;�[��n>�=d�SX���mDZW�8��d�2d��5e��W��p0�	s�nS<Q�z���`�\�m�H*;H�@���<4i��������w+��Jx������/�V����Vٹ�<��W��8呐�E�=w [�r\��i
W�sx�?�M�d]d�~�������Ց��f`�v��?�~x��_FO*�<����� ��z ��S���w�gH�kv�xt�Ry�����6ݖ���6Ԃy��:A�Uh�a��̝�J�#����ƶ��/�ncߎ)�=�\}���x��_��t���YYۘ�,�&k&��$w(��b��U&f	3T8�=�����m�;��l���H�:ü;�ݺ�������|��l������7�f�D�0̋��bnN#T�xf�U��t���zY�z�A��}|��<����ȭ�-�X� M��=/�0�XT�ٕ�s����k�K�nJ~�9�Z�~���l��l}>��nœ��.o6��c)¥����|�.�� kE�xxy�$bw&����..���l����~���Q��%B)_��#�Y] �+`�X�cz�r<_���&�g�����}���߮������af�Q������C���}yo��RQ����I[�wl����z�w�����9Na�z\~/o���.�"��uB���)*p҄[�>���Qs�ǒ��l=4����ջ�*}�ef�?n>�g:pr��o� �&��l%�;a���Ԩ�|�f�R��۷ѽd�R��Tg�:ܬ�|�(�bɶ��Ɲ�/�YF���Qt��.�iqNհ
t\�g�����;�j;9)��,U�KF"�$ɣz{�i	�! ����{����Hׁ�)�/���ۼZj��ϰ�^��w��:X�u}�!��^��^�r�#]�P����$��9]�M����;,��ۺ~h�zY����(M/aoܙ4���dƗ� ��v�<�f��޽�*������Ԥ�?Ka��s;)t�~��)�����������R�g�I�g_cꮟ�T����ĭKN^��>�2�!�m-}���~��ܱ���o_H��m� ��
�SR{1���+�	?������	a~�ir�Y
�����t�'G��[����ʁ�'�Ѭi��v_}\x�k�X�>�p?í����q�_!���%�+K��͍5 �0L�
�F>nX��jF�Q^>���� �]��G��|~��m��(�+<%���|�������Y�\��51~&�c\��.������(&JB��g��᠃!]G�F�oF���_/b���+��ر1�>��>kA��-"��x��7xC��SC�+X��JI\�۩)�}��L?�����t��]��LC\�Z��)�j/))��_�fE���?-�
�9�
��K��̟Tuy_�oݢ/������:�MYdaXNg���&�bu�����4>�"��۠���si�ߩ�~����K%�+-�E?���>`y�����!���$M�ѷ���G����vO&Ur�����:]����'{¸-����d\���,�Zf6��pSe����Y�շk	C�9��ی���y��m�S�S<�S�mn^���W�e�X��n0��4�s�ȅHe/2׺�ie�����=7F`B�}�rL����ߍ����>����͡\t=cb�Eia�̅��/
��΃��X�W����1,5ҫ��R���#b==}F����jO�&|czss���+�q�ɨ�+u��!��g����8�)����N�o������;dr���EM17�:cL'IHp�}f�nU�{�{� ��Ul�9����+�������o�"Q qA�p��+:5��Vp0.������0�7+�W��'��%���	��Rߥ�̜���˓�Z���5�H!B��2.��]��S����
�"����鋮�zoK��~�6����d����U���zˊ{K#{P�K��^���*Y��EM����f۔Z2��.�g�K|"A������b��I��? #-@a��`Y��׷{��*?��?p��H�>��z��R����j��Ú��� Oz�`)�)��7���;x<I�}�[e��-��$B�7���f*m��/P���	�8:J�6�]���ij²ȳ�C!�|y��L�4p-4�4�IH� �����:~�#mDk��v 4*�Pc�|���
�a�D�Ϳ��{� ��qY����=}��|W�y��Q�����#�Ҭ���6�Q\Ыm�K�Ժ���.��:{��3`��|z��[:Z���)99�y�h����M���U���>=�E�)#!���'���m;/n4�"A���������Ǖ�����c�g��߅������q�=�	�r����,V|J'\d��Q"b��iR��S |�-.AP�0Gf��Ks��r��fk(�cw]
}*�ѯį1Œp�zX�TWd�>���C6]�
�l�����{E�<�3|Ak�&�-U�=�5l_��\`�6��Ħ{?.�M�@���LR�1���m�72/~^<���Z��d�>��.>G.��|�h,ͤ��'&�У�Q����H��m�ԇ給ù>7*R�G��:���4���2:^�r������3��Km&��T���ʼ�Cm��)
t�Ie�w`l��[���~�Z4|D1�G�R"T�D��u�ݻ�5�<�i���V�r��	��-f1ba�$c��y�ͮ�c1�
0�R"p#]n�>?צ�"�tT�J����&��ω��{~��ʾi��v"m;Æ�X]�/�]I��~Jz�[���E�J�:2Y��AN�z���F*]'��m���u�t��|g�7�ߥ�����o��oW���d�5��m�)���_���\ gTc��0[z)��xӥb	I��N��6�l?���>���m��LR�6��W;��~m���h��S=���|ne�X�'�x0�G�����H����"����B�̕�#��&;��1��j�+�7Vz�������.� ��5��1��7��~����Hv}�Л5m<D������aT?t�|E>B.�ņ����AA����3���ה~[oL���D���e� A�|$ӗ/{�oO�tR�.��O"������+x�6A���ֈ<��^
�B▖��x�?j����a*�p�J5GHzJaG8�^+n�rf��l�ϗ��#�n�������\�7):^��i�i%��VZx<x�*w[6e5���-����-9wgRB7��D�`�ǚ��Ⱥ"1�{:5�j�g��QR������Oې��OX���dR��������{����BOdŜǝ!�:U=��4ĺ؊�$P¿��r�cՍ�b�p�y\0j�ٯ�t5�����}tu˼�hJC�e�D~�Ƭ,yV!�u(i� ��/L�~�p���~EX-�*�\��u��Q>q?�Xa��EQ}�	%t~�O�vYS̈́�����A#����� �vT�"���Q�Z/�`������� y5Y)���N�|����D��+�k)l��ث��d[���,�Ş�S!��)������]O�HdzIcd�ҧ�/z�3$U�ue�ڠ�&����_�NJH.*�*o`�,�(5�؅�T��n:�!��G���X	?&��i�GUұ��W��N��������C�Kk)�#��\BB	��i_�?���,=��z�PL�����0��K{�(F�6AeC蝻_�B��o�V���"UE��t�7�7���b�\�E'<�\�{V�[�t�mEÍy��y�7���g�mRs:�q����o4`)�g<�b	�(��L��,Fʑ'���Y�p{;��MV@�nI&؁�*줲� ��MH���I�1���T���������3xӘ�.�̣_�9V���w���rBU�{�Z���z����,�7�;�l��Y�E�9%x (Հ�!dϧ1A�Z�,�@q������F�ه,�,l���k�u�3�B������N�홑E�a��WP���]b����*�I�w�	�pt�i��vY�&f~���<r�~�<������zxiÊv�m�2�F=0V�mo��.ť�{*U-�����d1|�ψ<���9���Ȝ��/�&�����_�KzO�3}���0������=�nQK"+,P��k8����&�|d
�m��S.���]�`*Khٛ�bs�H���j�-[p���^�>��*���a�)L�0��dЕD,�_t.YA�1C�K�K Hip]��=��r��N*H+��X�lF��7�
|�0�����|h�~�{ͷ!��MC�,�
���	8*�c�!QzN��*8��+Ю�W�^�ꆢ�nV��L
�rd
DeQ>�;0M�iq�k�×�B�B�@ �c0�� ��sS�s�bҶR�/r���@��h8{�e�Iҽbfj:m��э,�&�%��@�ь�3(���I��~�Ⱥ^�Á�;C�(1���^c�4���^���&xi��m��EG����9�)���)���7�ZPʙF�? /@п�2��4#ў\(i�dx��3�$C:�12��b#+s��L.��Q������&g�e)
���(�D�L�b"���c�s4 Q+̇U]�ѵɠ��	J��,I��_��d:x�3.S���XgD�) �QM�1�tL��8������K�pB"�ED�\{F����	�u��t����sBntp��`��2-8(,2} ��Z^�0.Bf�����y�\��)��ʕ�9sg'&��7�3��)���y  @ IDAT�&iz�j!�Q�0��Pq��6��9���[ܑ�A �h9b�1��lWg;�ԓ0�a�ƴ��d�.:h��T���xn#�U���w&����8r�ic��{�_7n8-��q8%�d�F�*�T�$;Ǯ\>x)y.�%�L�V�� fҮ��`Z�'���ZZ�|.m��٥>�#>0��0/���Y`��D��������ln�ݓ��Ta 77;fZ^W�&����<6DFL���;�C��X�"������y��C��[**�9��#ʶp	�0�� �A�xL�<�<!�:��*P�P�ԫd�L5�>���OYP�!Kil�My�9�N�
U���\Q~�r��n|_9tD�y_x|%C!�|a��:��7��D�ؽ��'��� _�e�@P�g<�e��$_��
;riE���"m�G_�η�79:�Y}�\�Ðzh�Fȥ�I���������y8ܟP��L4�F<׫mm�`���r��˽T��/w�ma��,s�LMAmLOѪ��/T���˅�B�h�|��#8CBЍ��!�"��tQɀ|>������&�\�Aa�a- ���$
�����vkY.G*�+����D�u�����e����]�\�OEE#���+�I��~I�RT�9#)$�+޻J�#���ѹ�����w3H X$
�h��(��b"�s؊��3ef��<xLpi�\Dk��H��Q��F�[\�'3&��������]�aUz)/�2l�@r<j��9������ਬ垡]���� Rq�q턡[n��2eY�o���(k8���L���	�����@�il�"��5������褡 ������:�z	���.-�/tݜlaC�`'F�XMEH�d(�����&ƧtG��1�ϫ��	�"��j"K�Oh
,%�i��,G���X�S�(�8�@a�s�9	3��	+�}����.���e��2#���s:ވA Z�38u\WD�����!~�q&�ɞ��U�-��!Ɯ�\�k
��l\?RXT�uO��O�;i��56�ǤR�,6��J�Z&��<�>]�%:TD���'��CX�E�wa��2a(  �^���'����tE��8�2���e���v:�g����W�p�b�-4����	�K%��@m]t�5�OZw05M�����F�a#e`Ql� ߩM�[ᥬ�3_�0�&��}͠UdV����(3��D�5iL!X�"����􉃨�OS�(W0Q�
ҥ�7�D1|RU�ڦ�~�WF���R�d�ŗ��Fɛ��=a�3��Te�SC>L	T�.��luΊ#x&r��<_��~��j�j!GjB0��UNH#bE0�MJ��9Px"u���Z��$�05	O�['��I	�_��
�	]�%��^:�������Ԕes�I���	1�G�Kb��Hb�H��o���[��iɔ>M$[��I���gG���V��,��*[4��'c(� ���,CD��S s��z7E����=/�I����.ܠ��/�Z�*T�?Qj��pɸp'�	�R~L]c��FIN�ٰ��[��d'�GD��ՠ�����6��C'S2f]R�K���Q4�{̺E����~��lavz|x��$��)�I5�m-N`)e��9�UV2��ɩ�m41es�Bms��K��ٮJÈ��_[�B����aI:�yY�2�#Xb9�YŃZ�<���~bJ,a�ވ&:x|�+}�9dѬ��X��G;U.N�MV��^�ԇ�&�O��3H)��M5	U�#�tkS`ƼK/#
7�b��3+`���lbj�e@'f�;�^[�:�H��D��A���r��VqqӦ�i5DNNZ*�Ŕ�'�bU�C�g�>=���y�ʆ�I/�	�����,bE��71D̄��ɩq�����ʆ��� �)I�D��/���ҍ`I�%mS �z]�H
�
�#�c����cm9��$��>���ПaS9l���̸ED�H��k�E0	��,Z��-S��������(Y����y�rD�0P�g4	�	C�${ ���dFp�+%w���~]��'��R'�+U��S��F1�2�� A�T��e�j�;�T	$U��/�s8��_ʵ �D�^���3������K���ٓ0 fX�$o����&˶ĩ��dQL�ftK�A�dJ���@Z)��*�/�o�qa�*E����UMJx��B!%k0]zb�$�����O���� �L�d���G��A��*�e�2c3cL��H���7�g� �E5F2V�`�(n�j�x0C�.#��M|�ϵ��咯��ڊ�ƢQ
��WD3�ZFu�P�{��S��p���6c'k�D� IB�Ne�g��4FJ�H�V�K�>Bh��[�+��o�\/\=S{X Y�N��pc�r�q�{\�+♘!����9������Za��eV� }�_�R�@T���NK�*&�r�R�/�@���5E�FO�R���|55�E
�1)Ȩ�2}�+�p��)gȤ��.Hxnm�������D�"�+_H��$�J�Y�X�����I"��X����x���E�)�K�\���$�>��ye<�� 0�g�L�B���"�[�H<���]�b1\MBhґI>!ͅ߀��ҩ2)�䁾��Bbr��p��|r�����Ā"��?�\/,d�X�ɰB2�U8�kM�/x�X��IB��%�x�ʕk�*rM|�L?#�$��>	~ˁbF��K������*���%�6�9�%~�|%�ă�;>v�'��T������M+!��\��O.H{��W䳄�^��#�,%S���[������� j�r}��V�"^�0�q��I0��:��t������מ�>�sd�{��Y*���0��|EP�Ra�֬�S�I�r��`���H�#n>�|�>�h4����H�7f�<7�^`8��]�LKu,��5�]��I!��8{w%�T���J��&�K`��E�2'�g�)��͈�h)>sHz�̂�\�}��-	S���p�Q�L�M̘H�s���a��,�) |oW��N*�|]��t�_� d�Ik�F|w�|l¥�$Sb�5��k<-�(g�~�i�f�0蟚��=thxP�(��y�p1�o�h��eD�ܳuD3�\^�p���QϤ/�٫��z����9�6?}l�K�S5?���@F��˿��8�$�*_��U�p��ϵ1¥�f���J`K���:�n�;�
��x=��R'F,�0S�sܘi,�|u5�Ԁ���&�e�e�-5��0��̄��1�!��{�L��w���� ��R:s�iX?}��х���=Ku^5ts���үz *S�CDӭ������� up�D78�.�q!A
�L7�rCnBo����4�V 9loY%��y�a�����+?�^1�e�3�yK��<&���<�%R��<I�
\��,u	N�_����I	R��&���L?�e�6��+�m��Z5tSc�U�*�~�RqRRY���:�٤����e�L"N�$�Iv��JՌ��1�99�hI,K�"JH��)�6r�����P-˧@�10 c*M��X���i&vpBR�ҧ;uY���\"k)�KbY
��*g�_�63� �dP��ĥ�'��y�h)E����^�a�k2ҰG�-�aZP�!�1��Эb��\K�	U���$���t�Cl�n���t�3�������+��Z wȀ?�Fd�$�D��jMq�)tz�gr4&qM�G�����U����W��ʉ��b)������
��!�\|"*E�!q���{�_$0T_�JR����X��Q�e�bؾ�Ȯ�zٞ��r.��ϧ1��ӻ!������_08R�1�3��Bk�iX%�*ӗ1o,��]��:�G �f0!�!,]���Mf��@r ���BV��@<~�Q|c�+C,=��� �M��D�R�T-�>���zǝ����t!����{{���c�F�C�f�A��rsp�Yx�q%��A�U!q�F�=&���m�1|�%-7��y�1%q�����+��K<#q�x�'�р�"?�rf�m,�(�I�Sd<ү m���CQD�����T�\��O���=����8^�lݕh6�! �E$¯�������W��=a �n�{�&����5�x)w2� ,�G���)~up����+Hbĥ4�8��������?/x��g!�̨�g	�@a_�h}LP��)�牢#�K�*��Ew�EX�i��V�[-��2H��M�M,b0)�!�i� �2	�Hr�D$	J�z)��ra],۳���2�Z���~Źz��\囥�pe,D��}c����4�&V>�6XsKX��p�p�i��	��Q��%��^���/S�S��t0`-`��?��n5�1�QPzF��D��J&�o1�Y�ǒ�F��p�)��Ȩ����}���g`T�3�T;��T��@U`5=�N>��լׂ�v�,�yS��Z	�~t/�n�}w��h�!VU�;v���J(
X�b�F�E�S��8�ڿ9w�u�-.�ֈ���I���%a�~P?!P�cN�Tw���}�e��})��	�V�]��LKK;��쌃�������^23?2�0�c�[��m���ZԴ{�)6k�;��4��M�X�E���@_oc]�{�����?�S?���-��vJ1ri���\�D����2S��'t���Fr���|���_,,�8C����������ӷ��-C������S<V�g&�IW��A��6���LM�š��u�z17�P[m�,{�;$��bynfbj|�կ|�?����_��ΞMV��s�����,����!m��)`����KeU�AD��Q61-ۚ�X�85>��H�ʕɑ�_������H�e��s5���A���A�qx�q���\b�m�bm� {!��a'��/����=���w��?��-��ih�����H�����1��������QW�K:f�w�;���K��e/[�|��������~�ۜϰ0?��I�bw�
ۂ��L�IV���
�&]�^���F&����Nuu4�����{�}�[��ƚ�剱A�,�aCVb\6j�&e��XWo�P�Lg�`Vt]�9��{y||`~~���y��g��wݹ}�f��5�-��aav޶(q�hZ�Ji9���%�V!Z0=�,S��F�i���ZRΪ�ٕ����m������xe��x�c�bYi,B��[�\U)��՝��x�&�ڏ�%�E.���*���zzft��-���6|N\�R�&'_�=I�$�	�a�W��?.&�Zi/�P2!ev߱s�Ѥ��}�\sÍ72 �;fs=�G��,�_I�d8�K+��h�<u��ӂm)��:66\r���u��{�O��-o~ө�����^sͩS�N�<&m'c'𹡩-��(��K��Qt�;�Cv�=Ԋr���6���/����S�'���wغ����6Pv�g��yɦ�689s����}�A��6����2g`�=s��]�WW]����������n����[�F�\��ơ�eᵷAGg���s�����d���im�m�G�����r�ȳN�����߾�u��}�m�9�xtl\e�+���F{�v�i�j�M"3z��~���N�&*�����_���~���Ů�6���~�km[��Ï�G[I@# NX d�L��ʢ�E1��p����`WW��cc��������/�=w��/�i�U�|�	%ڒɉI����5	�nβ��p� ��ο�յ�L�1��P�e�~�#=[6��7���
���|}g��f�!��� 3Se{�rQ;Gx9*)�*[aؙ��x�/��/L�����W��e/}��'���wDD�1ئ͛�;�'d� . I\���+ؾ}k��:n��G���:(���~��x������?�a��������!<O�'��%[� e��b+?1��m�:hc�������o����?���]�`X��CړDi�َ��_�5�����61��l��Ρ��u7\�̸zGV׎�9������[�z����5jQ!|,˗������� � )�W��{�n �9C�iG�o����;���>|����8�a�f�5~�q��ím��c ����s��!,���Rb������eO>��\��h�H{��=��O��Š���m5�չ��/|��+gN��������7����>6	SA�D����ֶ�z��ǿc��l����;����=�c[���pCckC}���s_���-�pT�,���7=��wEL���m��뮹~r|���36x��������S��~�#�iji�ٱ��|������E��+��#L|9t�Y�J3�bB�i\۵��l9x�pKs{����8v�����}�����������Fߺ���}��Ɔ6S5b����/}v́�I�X������c�ES522�窝���ںu��ӧ4gf��=S��ۿ�{�܆�ͽ�g�l�1�ճ�Ȃ�W��L-t�5�\s��1(�����=��|��>`S|G��tĎ���t�ׇ?���o[�g����é���{�'q>b1xqA��c�}�}���^SUg��:��}�{�^���Ǐw����݃�#���=��w-p2a���vD/���{�q/8jD�s��S���o?x����`��!%K�M���_��3�Ϝ>i�Ʃ�'=��߸�a����6��h��~���h�R �t����/}�;�1���,�򪗿�=o?s�c"˖g7v����9���2�>��[B�+���іj�S�,&�ű�Wm�������}�O��rdu��"?UZQpQ=J�Re{'�.V�ɢ��,z��w�\�j���;>6>aSi;3�ʡ/�(kQ�DfV�P9*���;x��3Nn~��8e�6��g������;�g��8;�Lj�캪�6s�,�[�h?=Ӣ�x"d����ɓ'�@�ӳ��@c[�?������N�+�t�K��]Z�ؔ1,��K�b��Lϵ9	f|JE�-{�UW�=w�'�|ի^�m�;�,�8p��ѣ>��'N@���M�ϞQ?*���W.�ت��;7�E#�o��x�CkcA����8ppddl|,�_�x�0��7�֊�����9wH�'L��|���[�DE��uy�7�y?mEVΝ��B'O��n`wE��j�1��I\5�2�9��Q\|��'���Z[�Q@u�M�8���{N�9��ɯcG����n��m�t�#�!�Tm�%���g�TԴ���}���k�ޫ&FG�;w��1�ȉ��p��Q�6�0md��ޅRilfge��|�d��L�����7��]ݛo������O(U>���gY�9�e�����bn�LOC�����w������K�;w�!�q�<o3BO��>q��C=+��ηa����D'_Qjfm�S�}�v���ho��@������s��%�hӼ��!�%���=W�ґ6�c���#��e�č�=��c�뮻�[�T�O�����S��IeT���!9�,����d	`Vm�sl`�O���@�I�<���}���>���ͳg�b���ݒ9/Ó'O����c�%��f��K<�����Iȟz��tC�Nom÷x��~�7~�Q.�����;~4G�a�X������c�G�BT��w��ni��[{ZZ[����ݯ��u"�����a�����+��8����S؎s��IZZZ�`6%����iu���X'#]{�5�'�x���>�	�pˇ>�j������W������F5��C:}�|�_�*��ݻ�y'��'?�����`�G�N�� ���'Û	���BfN��9`�֙p^ၣ�?��[{�9Q��{�����o������~�	��<-ͭc���O����� N�L�~��s9!bhؾDUwx��G����[{z`�K_�k<����!'}S�=���~`�~��.�X8�W�'{��3#���b}(R��/��S~�w?z�=}��	�$�>�Uj�C���{�D�y+~��6||�h+�C��?���ww�ܚ�̫%0op`px(�I��2�c���|[���hWw'g
i�?��/�����'�<p��72B�3Z��ؚ���Jj��~��1gRb��9ml�����Ax��ѧ�|r�������/�hǮ�*�jHJ,�l��a����� B=��޽��E�h�v[]n޴���׾��G��ݿ��p(C{['^W$^(}����9,;��	(P����8a\�s��\0Y0�|�o���G������۱s����Q^�!Y	���%b���s�
�8�r�Ƚ�;��������=U�P�я����~�V�M�ӌtv:[V����a��9�����q�h���x��]ΆG}�A@�{O��o�W�
��lsh4!�tA&�d)2U?:,xKQ%��<įՂ���v1}���]�v���}D[����z��@M;����1� ��B
�)�G�i��3��((������>����t�w��E~�w4��^�@���+O�$_u4P���k�V��\���������/~k���s�	E$���Cud�s�n�~aC�5� ��5���ͥ�� �bRm����;��o2Z[ۙ�_��}���j&��jP�-[���6|���'F޺���2�	?0ĨW���W�&���^��'8�?8�?��Ƅ�9u�/�Ѕ�dަVUf^�&�ґv�Q����p��jn��^-���䧀2y�vf�sA�|��5��C�Z�>�}]E���G?���>���fؼ��p���kC8�V��O(��6�M��/T��f���&G��s�W{���If��C��ڎ?r�X8?O8$��WŏahŸ�����C�ZV==9u��t�������t�D��mnk����з��v��>TT1��a^����F�G&���hhl>�{���x����:68���<�:�s�N4�����! \�q��vTl�몋Q����7�y���5�qhX��	P��g�d�'�z�#U_566�x�Ʌ�980r�����ttt�;�O�ٖ�O<��7^�L��D��a������w'��&Ua�{��w����=�����2,(D� 3*hDq�	.Q��h��<�$����$� �c ,��1
��� �O/������;�������=�,�<S����[u�ԩsN���}O�ݻw�-��}&U�i�V���M`���e������vGʄ������x�y*6���V�	�}��Q%���3��tF���M�]#m��L��x7>W:�]}�m��pGؗ��t���N���2��o��'�n��Sf-R��u_]}$;��F���̟�v������qI3<���/�����1@����_�º�.�b!�͵L�*�^;���&t��]�S{Y���F��
[H�?���!)TF2s0��x�2�NC���gH�@j��Tup��:�Ԟ���V+K�X�ΝϺ��r��5�҂���'BtR֝k��a��FQ�i�����o�Af:�!l��z��oАǌ��'����ʉd|���֟@>��i2��&�ٳ|���(Ǵ�Y�i�f���"��Lh��x'Qd�!�T+t
����9��N4�R���G��6�Š�Nh|֤�H:�q��M�q�т� ֺF�<��֭�f�JlZ���Z�P�Z��3���AV*;˸�?p�|B�h@�$MŬ%+	-??��x�̹�~��L�3����:�rյ�+o�F�2�?m��Q.m"I�G������;�Jk�EH���+ytݺm'��H9���0���D.+�v�3m���M,4�oUe��KV�qR�
�!�)���D�J�BBs�7_O��P�J���;�^T�_B+!o2�\eB~�O�gN���#���QF	�ֳ�)+��5l�6���:�
̂B h)"j��4�]��)5��:u2��E��K5ac)�Cf<͑6��0:�G��0 ��9$Ю�d3h���ή����.�?8`]�C�٨���U�,`�7��Aw��i���.��5!�o��r���)���"E�n�@����.8c7�'���q�|�ރ��>VF�x �h�����b��v>�)�Tf,��:Ϊ���lē6̱�՝�3gϢS�L��I�ݷ\�p�����3�a��{M'z9m�G��pV��E�U��Ul�{n�L�~�cpu�#���<gٙ��ԩ=�
3g����}���YHc��ԋ8�H��ᆅ.59[��*��XK��,q�SN�B>�?n��+B��)u]��ZU��\�)o0�0*&I�ĎI��Ia�)� ��j��F,�.���έ���[^�3��tې���F�!�A1+B@W����p�(�|�[3\�)Hc�l7���t^*U�����*�]��+T��!��.U'6n��[�����D� �_!��-|e�삢��y�&�hɐa�N�+�>̄֌~k��0��U�*lZ��������|hz�x�� ��H01��>�5p���|��_VgȐ=ƫ�>�i�u�O�B��3�^I��&��ף�Z��b5Z�n�c�[i�9���5�R���HgH��!;�u�e;�P�����c��J��F�ٸ�'H�𽓑�E���e��\2�fo�GI���u�ۋ�`^��fl�H3�g#:%(Zs3Z��W���/n �$�_�Q��8
D{9V�NB+z�ů<Q����-�2۴ĕ c*�t3ᇴ�/B5Z%�P�@;W���q�@rǠ�8��T�
�e�N�OV���!0��$I��]�ܻ�nHv�\iɦ�JM�ٝ��>��f֒�����/��p��)�H	l[i�4Y QO/���Lb
�½�AOh4
EbX��0꺃�mDg{�T��ID�AeZ���\���1�����/��=`J��G�2E�"�n%�b7���6�`�L�Z�8I¨V�oq����{���lf��1ZѴ�%�ǭ,�C�J�p6*W�.eԝ@�m:�e�N�+�5j��N5l��� ��i�_�1
����Ș����v6���Mb�<��$C&��2$a��`��x�݇	U,b=q�v,.���X��k%\b��YbT�K�:b�2;O�,��i�)�u��`5ڊhA����8K��V��ǰ�s��c���袢E�*�d��q���]��t]�"r[&�K�Ze;�Iox^k�56:�/	�4�Z�.������j���Wʠ�D茽{@Fc�cU4�ᆒ���Q���\�s�!Щ�!jD��� �M�u�������{JP�*5��	!�}��
����h�XK۾6�>$'h�r.��R'B��/�$Fat��q/:�F��rԎɜ�ٽ�k6�ÂM܈d��d�B���z����r�r������ ���u[������v�M�;7��ov9��!AB��l�Hj��i�D8��Z��o��K�K��x�-�{1����i
�h�p_T+r/����� X�P��~#+�y��ߩ���TR��HHOy�������	��uB�S'�
���5�S��p�l%ʔ��Yf���TVNjtn�Ż�9Ń�T�aA�����a̠�#�U����	���d�(�T��m�*^D�cHr��v&A�U�jR�j���h'ԍ�ak.kO�m.�C�԰���X�مl���[����:1ށ|��ю��	$괉���2����Tvn�b�"��6�slb[��Н�.��ql����� D�U��e��b��IE���MW��O���������b0UGU��*Ӗ�b�zh�4$/�^�:8�\1��݁|Q"[ǥ8Ç>6=\1�f)1�~ghF���UNYS�SfXN;9	'/����uE���sΥ�G�l'R��l��\���Y��\,�9��7vORػHQ<^ջ�e,gIF�y {�!���Fb���C��.��[�[�Q.��/&8���'�$���o�B���	c���i˳2�C9L.X���Z|�����R|���e~�e�';�]_�$�%�N��7�q�p��fW���X�#C� ruJ��]�mAЄ��f^iB�����T�V\�Jk7z�E�+ь5�篭��I,�'�[�y`!V��҆�uO�M"�6t���ۏc�SdZX����
���I�j%r23񯼨���T�Y��!�#4��(i���d��(�'��2�=�=e�t�<yI�Z�����J<��F�`5��g����y�u$�|,�Ɇ	��Q%��v<f�W�	��i��b�R΄��*����
>,��Z�ΉO�:�Ya��f����x;%��4�,nmI�<�	����'w��R❾x�}
�_7��yU�'���$I[	E��O�
m�����	��#��=��eVO�]ho��^Kh �?uѱ.1_��/����>Ǉ>g�_��i��G`Ҡ��iw��Q��O�B�e�������GO��N�&�nTl�"md��'�����ڋ����9�Z�x��ꁱ��
�����~�{�q��iS&��;q��]���Xeς��s�`�X��/ډ�py��c�<@��sVnʊ�HA�+���)�����%V�-�HO��OE�Ez
��B�����s���ԙ3�l�������0�$��A�މ��p��t&��E��_���b�41�ǰ�X�,�+�%�1�F��I	��b
��o���t6�m�~��A����&�&��|C+��ؖ �F�8��@l�|!!N��iL���d�$���ㅺ�ԹЏ��Z�z��*�r�ߞ:ہE�H�i��L�o�I�Q�)�����\`J7>m:�]:��.�������B�
TEu�筸[W�"�P<C�s���S9!x����VN3y�,��]�x�$?2��0�65j����%����!4W]�NW� ���:9��N�ЉmNxC�t�=o}�/9Zs� QA1���t7���P+�hv����E+�&�D&�Q<�o8�=��Z�X(�Y;2]�������uU��w���P%��-�iĲ�r��o,��95R�5J1���EI��F�:HG櫉����"��pf �yU��S	usЯ
��
�Hu��V���:��p9�]��S	_��fJp3�P�����ae�b�v6�]u�*�_��-���u1�D�j����C#ZJn����RB�b�4}H�˸���w�p6�+M������k�E"�Q]���d�\YM*9��8i��7�nr�z(��@S3�n�h��V;Cy��ZPU%�%DpI�x �%�USl�h"�QC�j��$p���{���Vu�,��f컪���BW�A��	��'����8�K�fՂ��[P��Ձ��m�L��t���V���\UK�0E���Ɩ�Q��c�5�h���&oa�)�P�����h��5e+�� V�)^�6�L��]r�NT!�9���x�G��cv�v��;;���昣�M��S�1vt�ū�d���0@5?2�Y��a�qԷ�lQ���@=� ���#-4��A5��� �_��"#�ҥq�-�8�d��~	�*Q �2����h���ZjhS�v���5����Ů$т���T�����Se��Xepa��ߥC�� p�Rc�	�*�1�f�E�B8cc?v@	ۘc��R�96'��@����0%#fo2'�vBTay�͙}�h����Isuc3��������ٰO�L�BLL�!^�v���h.y1�^ɜl&YT�㢩��BR�{Q=�B��6�H�)zY����y2�ouUڑ��[-XMP6�Y��D���ܨ�����\[�L��+�tܾI��+p��ty!F4Gv.�W*��#�*�M1��N�nh�LS5�". �'���l�) ]�v�ꥀtz�v��.��z�	��m�Ǜ	B��@�yc�C����] ]GV�t�+Y��jW)�0�dT"� ���h6���j%jՄ��#��+/�v+�tbRW�q���d{���Jd����h�N�Np͔�;.Mw��U��E*�kb����o�&Nu��$;����t>T�t가�p�b�(e�:?�S֥u��Qe)4j��h�
I��
ը|uj�]��*�4����p�JQ�B[�	���~��e��U�WH�i���]�V��}y8�����E@Gf4M�و�?<�)��SXcƐ�*��I���&3�)t�W����:877��R��ӕߌo�!ė4bK6����ع��Ɋ�+��6�[\]�:
H�h�ʊY<�HF[3�Sp�
\������3dI��=f��ZZ'm �)�l�|�D�!6u�l��[�7�u~b�5�1�B&p��u�L�� 2�Z�����TA��U���ho���R�ﶵ:eƀܹ���c6��4V�S@��0} 7:�ŜP
��h%���!�9�r����j\&�c����.T��q�J��D��WΕh/�X�M�@�뀪�-�ʏK,w6
�,.�]�|��sn�RjDh��BE�,$�˚%n �5�H�u�3�O�b�X�e3x|!�N7"ݣ��9l�2!�m��%o�&��sU�z�=���`n�8���ӯ�|a��G)�ޚ���z��i� q�b��PrIإ5&A{A�{'L_#�@��Cg͜�1o��ۘ�x���AY|pL�uXA¥L�D[.�m��2u
�F��<ʜ?r� \��ڵ�(�8�Ay�A,90|ԇHh��ؠ�=���@&�]��N����p�WO�iq�F),&�|�ק�>���u9��z��Sω��3L���'q����)���嫰��х�s\UP�^d6�":]_��u�>t,��$E�	P��.���(�CM p\0W4��ZG��u�rt$���CuL$��ꉾ=�<�z��:��H�V�$[ɺ�Z�,TB�����M�/����eO�L�eq|mv��#xrN�A���T��	�
@Ưd�w-(Yl������1hs6PҮ~;��V�I��.p��s�Κ5�|bPtLJ僫z�6���:�NU�>���hf�=��-9$�$���c�ʫ��6�Ϝ1�k��Ǐ��Vj[�38��(������͜9}�^.Ÿ\�5��P4��VD��M���N�'��Pt�;�r�0k�����g��U蛬O��D�0�$����	ԁ_QŻ�}}=~�J�k��"t�%:��{ ���N��i�j�|���rv���똷;Hn��lḢK����e�y-��lx��'(�����9��m�nhE�b8��Iy����y�(�b�x�C�$�,�LuM"��W<)�TJ@Ę����Ù�ah���у��ŗO�����s������Фji"X4d���h��!�߁��a�����!L��"(� �@�z�o\��)�'J�*
� hU�n_���}#]�:fw;Q�hs���ho.\؁ǧ��d`���ٟ���Șsd"D����'W�]����h2�3�;�/������yJ�@/��f$�Ż`4=��NN�*޼9������㓗\�Duhh�Q��>��!��#!�dƌ�|dU�Pl���
�wK.�o̞ܴ���O$ @�=�����z����,ǹG�<r�6�N�����W,5*T�5u`8�j��������$�W�[/�������O]̼���( .+�T��6�ޭG���i8��˅
cG�O��m��"�o	~[����]b\�L|A>{�O�=7h��t�� fV4mb�����$Ub\8�W� ��G_����)G(�!��}X�����6�./���W�Z�=g�߿�|hb�={wH�+11�����{o-��0�4� �<���x�>(����0��^p���"Z7�
̘��k�)و#���1��
�Tv,ʇd�3�x�	&{�J�(�0�a����;�����[fB21<�O�J����ם�[�/>r���@�ҥQ��	��x�=m��)T�9*Ɔ[��l-h�.=�*��!*LM��üdsҎ� {@��=v�o3ӱ�{�����e^�a�\LS"!t̊�=tR��x|h���C�9�<u��ߓO��,���=!��j ~��-d���㛁Ѕ	��RpzM��������$V��$Tc�Bð2�fF"]�nX�ۂ�5��^*�cit�쩂iǤ��z7�2����=� NB�����wΛ�w�S�b�f����f(��9�$iG`y�6  @ IDAT�2w���Mh��W��u���S��L[�x��f��Q���q��Չ�l�;�v�P����?��v��B���f՘����l�, ��L;���R Qu?���c�z���B���"-t�Z�`\�+������`˖�h��-�4`�±-�
������)K�2hi=.�9�[�|�_��g?�6̺c��ѓ'��ݳ�rTm�`���섺��g6Ϙѿ~�c��׼����~����S'�Z���y���l��w�G�V:�����{$��+ҡ�w��}�W,~�^{�sn#��0l&m�*z9�&IL�D�����:E8�!3'�ݾc�/~��������\��?�H�)c�ꦜNO�&>.�8�������߻o��^�7��{M�;vn[�hh����x�0����o���Y�f��7i��];v�޹��k_����g�:{�Lk�C�jS&D7�:� �s�կ����i�3����y��o���U�y�8}��R���WeV^�.�=�`�\����ܻw��y�^��o����hZ�'7�3d�R��O\+��4�٦�pl@�����z{'ؿ�N�-7�}�n�� ��G)]1�����u4F0����ԅ��̴�n�iժUh�_ ��Jb!	��x�k�Ӌ��O�3�{��͞=��o����鼪��ya��}VI� <�P�/[���U@M�) �gȨY�.Z�X1����g&O${�/x���ϸm͚U0۸q�6�Ϝ%�����c��a`c�)�ؑ�C}�?��7��$����G�?��r�ݯY�dэ7^�u�V��Љ��>3g�<�q�'���0W40a(FD�n�R{v�%����-X0���׮�~���l��*�w��>��!V+_$m��٬ Cbj�1ih�U�~��^w��7�p�7:���͛7���P�L�x�b1
�Vn�ls�5��;)@ֻb^˦2L�o{ۏ}۷�������{���B���_p ��³d�.� �ŜJ�ٳ��f�P_)|��^�X�k�]����(���e`r�6�Y}���&U��5L,ޒ�*Y"�ж��;������/}��M�^ö���os7
Po|�<�t�R����,�B���X�>�TF�*x���"�Y�v��|���Uw�^s��Onzr�.�_p&)0��-�'�]`��]�h��9ad�D;�.�������׼��[�tъK�ڶw�A^�
�P2Hg�GR�M�A^fW�{����'��M��\���o~ӭ��<8�{�������@�g��8�AH���ūx-���;V��;29}���ߴ|��M����MM��;���in�{!^�il4��`������=t�^��w޲jӦ-CC�o�����{��v��=���;+<Tϴi� ��S��Y�b9:j(��i�O[�`�[�_���t���gܸ|�5�Ǿ���@���9�Z�`Q�{<���0S�"���ќ ����e����.\�9u��[�z���{�n[�r{A1pt�J0�����&$�qe��?�=��~��0��Hy���?�yw�V�aXy�A�p�mi
E��B2���}s�����р�P��׬����=�9���Y��n^�l�qs���t���&��˗�Y�d¶�%���L�U��A����W��}�����X�zՂ�j��E�����(�Z�Ν����;(Z��X�zu�y���d�$^y����'��������qn�W�_�l��ݖ'�1����H��]6Fpf����}��-6-ں���t�w���oۼe���7ܰ|�r:�r�H��ځ���+�S�����:Уנj��c�uf�讻^���˖��-�-_��o�&'.����a�6d�7S�a�t�`r�̞�A=$cp�������yͫ�����̞�у�N�����%��B�M���G=����|��9n���q~��O<18}������W�����[	J�SЂ�E{���h��^���b̈����[�.Z������f���o��o\����/_���G]�x�K^�'7ny��/� ;�p��9q�R��ŵ����xɒ%�?^i��衾;^��o۰a��f��~��|�-\(nۊ���M�K��fs�͉7�'����i58Q<J�H�KMk{=��5�����o�|��w�񒿼�S��Hf=�Y�x	�<N*$C��6K�,�I�f9뀝;��r�m���W�l-7{�|�*�fc/�aZ �؈|jb.7H���2���z� �p
K�.\8t�Mk/Zr��a^����_�+_������q�U�������x
�z(�uXk�FU5^g'�g���O��o�6��?���yC��X�r%z;z��7L��q��#-r|Gv�/� �ƛ:�Ю]��Q�;8�=s�曯{��P����=�����g-޳��_��h�#E�OA��?�$��ql����!	��X��/~��w��ݧp��m��_��%/~��?x��1��N=�h$iՕ�٘�&91\i##�r���_�C�:��v��f͚�A��)���]߽{�S5�d��~9pH�=J��`��Z䥰�.Yl[����F ���<�2�����9{:lf�#�v�{��z*�_ �+8$�j�a���`��.`I���]{&N��z�u���������z���s��7lf˙��n'��5Ռ���wnݱcYd�ߴe�|�~ի�����M�׬�������/�?�����C����
,���{�ETB�+����Lڢ~�}�����/��/����V����~����cS%O��c4:s���[�l����2I���|P�h;�)�̞�[�|͝��3���C�7o����?}�c����k�&��a◾� �ࠉ��Ə������nk�q���_���?�3?�f�j6����?��O������GQ��M�ˇ~2�I��7⳧M�文zH����?��{�|��moy˛�c=q����[��ǌ��3q��zd9�D��v��=1��`Q�666n�h�1<�C�G�G�G~��/~�k�]���|�������%ޛ����F����������P�@Zpl��Z������L��;�<��������.��p�����y������b{W� ��[��6��[����my�fKJMh�=F٦M��{��;;i��5�>��w~���~���Oٷ�0��i��Ι3oÆ�#d��-���t>�|�*f��'�x�֙F؃��۶���o�喛������ٟ�W8I�Z"�mg��u��cx
��H�N�1=~��"���uJ���xb�x~�-߷p�����!`J����2���.��t�]w�3[��s!�9�.X���mf������{��뾾�t�"6E�U�W9ڌl���[	�.�Y>,���:��PاO�.�9��m|ֳ���O�����{>���H�dyC2�ܜ&{�Ŏ�_�mb�D�A��Cx���cs~�K���������x���c�a�C*F]Z0D��Ti��D;�Hʵ���%3$���#`>�У�������}�9�P�*�הEm�F�Xki:�e�ec �M��Epg����~:,X��}�������������ʀA��ӷ2p��?��Z������w��?��7�488�W~�ߓOk�-[�͚9a�لo�LF������OσF1�e%BM�w�uk?��O|��������$��aN=ѵ�I�9d1(f�U+W�eR5Z4 6���O\{�Z���o��>�!�eHB*pK�f][�}�q��a$ŝ�Z�?�~�tv�@���n�v�}_|����G>�x������0�9s�Gsz)�1l+_��-AN'��q���FjY&��XA~�\�z���չ[*a*�	���6.�!C&ю�4��+n���&g/�����^�ڵ���=�PZ04�%�ǾUɁ}�ζ�% ��@�_ 4N�i
{��Āg`G���_}�.òeC>@��Wj�!���2q�'�P�@L�	�̓	�9p��uD�#�(����s�O�Ԫ*�ڢ�U3�v�&W׬�u��o��Z��[o����}"1�/{�.\��C�q,��0*A���S J�����>�u���|��6~t<��^B5겻	����
TG�}� ������Id�0�D�~��ҍa�m�n�m&����~�r!��'��x��WpT�Z��t�*��c!�x"��#�Q��|شi�|�2q=���L٪X�Ŕ.u!��� �Ȯ� ���'OZ�lŧ?�F�U"�B�����W�6e�8�%%���0F�V�Ja�֍Sm�g߾��A't��/��-;��,�Ȍy��y�`,�;626l������)_����]�w��}Zb	TQ�;�:��8��P�����?��S��v��byS�}
�U%E	+t�PY�f��3ƌ��{?�q���U�{zb[���7�c��F������P�����+(b��ņ������!��F�c(䨠!(�V�!Mt��Z�b�-&�d֢)�D.�T���(Ƞ��%(Ώ`�����y�GIE sS�c�����
��
ICE�����S�~ E��%�e��جY�����y<!���p(8�ҝ��3�E(⸥#��|˖-�o��<4���q4}��*�Q4*�-���xi��;b��4�P�8ФvG����I���@nC!��@)z�	n�	K��86���>�5/D���?�`���^h�.�$,0Z� k��O)��Ei`�h�&���������y �  ���:�ML�>�J�TG�1g�Z����7�1"VI�_A�e˯9q"@2�v��.%j��fY
���A	gOx��;$f۶[�n�c[1A�LX��M�,�Ew�l�s��Q;��M��V��a�D��&Ȳ��/;�^U:��A�6�ުH�p�V����e��H���Qud(��C��E������v�jW�`䠑q��||I�I��YkB����j��Siq7�JW�"�Ҥ�&ຌ9�%ӥ*��[��.;3���ۗ��,9��9�8�%��P�1* -V#a6Զ�0���)F������_s�5'�;@p=r��(���,���0u/]L����)Ǩ���.�̙�-ؖ9�ŤmƋ�D��3������b�!�3g�u0���ѣp?k�ǽ�P�m������p�p��f#�O��?�,;>Mg,�K���v&�b`�*�F���TU^��zHD�crUp��ƥ�!_�8ыSv@��tjX����X3�,D2\�����ڴT�5#HG�"�e�C���B�]�O����f�]�<�G��V�W{�euZ�:i����X�Rp�N�.���\ZaDD8� mi�떻Z(�m�R�!f���(������Jb6����;�ʝ�Q�}E�C�K3��"�:j�G!Y��2��qmIԸ�4^��J�esزܳ/��'���B1D�E�����av:�б��9�e;OĒm��n��V�~*e�����GI�1LZԺ�,���g{�Λ�@[�D���k9F����?c�G2c�Xp�/17��j�J;�q�.zMW��?���X@�NP�$�nR]�.���*!��P����m����<]Ol�y���3kb]t�=S5A3M?�b�^�-���.T�4H�/H��:�(-eLP	�J#�$��8FsT ]��~VZC���6dG�+4�A����2Ҁ�(��,P���+�N�*��q��v�.H�g�Y�7@��Q��Z���lU��Oٙ�� ����]|�P��5��v
I۷�c��>Tv�Yf�Cu��	gu+h�eK�*ಂ=����-\24��e�`�|������
 �8��V���{��A����;6��zɂЕBI��m�8~�╬0<�Q����d�~>�;h��&��濇�t�����]�I��О楁2�^d���Q��>VB!���.Y�`�{<C,m�Ѡ�Sev�_�2B�|!𰁖1�m�أf�fC��d@_�y�`m�j�;6�P�@���#�n݊#��b}&l��u)n+�J@#ȑ��,U*_�֌W��X[}T�.�nw[��O�ȿ���,.k��^:���\Ih� �*4t�0>�a��B�e崷چ�?�GM1�z��	ν=p�gWs��s�"��>�c�*0h��Yޝ
����0���5�\��hK3�؀�$�]�*���^v`4�X}D1�������u��g��rxD±��5�;�h�\��I���d��.�m�p/�[��B��\���t@�p�4�N�	Prj]�� 	2�������
!<@(�* ��2lR2Iw< �]5�;l8_5(~VŐ퀻�׹3���~25FQ+��Մ��|ERY���bF��qV�!A~Hف����&O'E�tU���"�NuU��	�kTE0T���x�+�Ж��4�`*I���ŝ�qY�HT�*����"By�@x�88H� lD�ₖ]����b&=#��م3�%�7�
��Ms�o�2���1����-#u����;Њ���b�ɬ)v��j�;1����8ZO<c��N��x�!cJ���4�j\#�λ1�
��D](@�#��X�J@L��O}���x��0/������g�gTO�V���p�]?��EД��q�a����Ԣ�ܪ�ETO���[+@9%8x��!�&�'�={��m4���q���/����F?ti��V��73�9IͲjL�-�i��D/��� �?m�(;v�X��Ӊ�(аG���Y�:�m)�$�r�<Z)Ǩ�!S���u����i��b�,�1o&S�Ã�7f�6sX$ڬ�$�D�]�n�P�x�*�T|�G)�'��J�.�]?"R����G7�Mޫ�g4����&JFb�N�B���*J�	��Ŭb�MѢ�5��&F��3�.������:���pCu�t<�U��5@�1Lach�r���V�^�������Mb�_�#����+���6����O���#�Xp�g��b���2��Gk�X��!�����jn�Ƣ��J�!zE	C��,Z�YdWV����;�/+�V����)B˨��T�M�a��f�ع9�V'�鿗� r��U�Q�.���ԕ��A�N;.g��]���v+�ϻ#��]*��;mZ"^H��ct��_�Y=��M��Ȍ;�:� [m�`C"t���Q�]G� �Ӣ@��Eގ�L��*�gܪ�L�!���U87ǬK�G:��c���e(��e'{��Q�O_�=P ��Ď�?�r�h�D��#[iQ~e˧V��]If�%9�4�ܕ��������R�>j|[Kh�c���H�yi(T���4�U+Cp
V�^���S���U.�hơ<;(Ĩ���j*FVɧ;׭�[p�����ET��J��Qe�����!��d�l��X�]�'��-�(���9���<f�Z�P8ӣ%�L��<���u+��2�N�YրO^���B�mӯh2:r%ү����F�h(nC���ʬ��/P:q7
-�!�Y&���O����4�c��ob���'��;#ԝ�t���,�8�$	�$6X9�	�%MhUy�����T��h��.pE@��w�¥S<�dٚh<�03��4ݱx�əa��W��++~���3��e%Z ��!5g�(�%%5�jձ��bH��s7('���ml eǍY���-�Ҽ�D=	�c�粓��A�1�G�W�@��B֫k��Khl�K�(�E�3O�S�F�rq� =*&.y�@����U�.[8u�d&m�&�}/�8�C�H� @��>6w�@` D����'�ñ{r�5���������������!��4�jz�v(�t��[�F��_�<������!����l�+
w�+��=�1y�/��<�`�a�^�=:-E�N���,@+�qT�뼼¨�"�ZH"Ep|/�]U#qx�O*/��"u6��$Ϝ���=��Q���gN������Ǽ���5sr�Khyo��#Ϛ����%"��.�w6eϨ�E�bdF���s�`	��4.�J�j�@g�Re���0`@` �"l���Ɋ�t��ʗ]?w��� ���sfL���6��^���9�aHg�y�i"�LE��%��*� EW#V �� ٕ�@���Jd,��	.���>���Z���,�%�t0�������zW�[� z
���|k(��������<ͱ��"�`Y��������g��.�\t*n!{�������_��o��̸�/��J'^ ,J��1���;�2=���[���r�&ȹ�I��<]3���^�?ط� �_1��`�8Nd�]�-���3�-&���$�cr�xx��K��Ɨ�ǨeWǌ��]�%$���J~�cT=�&s<�M:#miOf�hԼ��|Q_u<��"�KR�V不 (�,d>�V��Uc�:?���Q�, 3p������J�	�l�$�Ȇ���DY3��Y�J��]�3��$V)M�M���p:p���)�#���z�(��� ʤ��(�a�vw����F�~�ƨ�1^��
���q	@]v7
�S��VvN�:�'�M���Ja�/�7�SK��6���_*�KDeJ��&v�n�ͬ�U@�(`�G�
K������-RIBB�R{�Bsc�}w�P���6 d���33tk������To(ո�"�ۼь@�è8���U�&� ��3�4	,�Ȗ��n�`�T�5#
`nL\�FPF�hɦ���]�IP'��!����A�yi�On10���W@�3�u���.GR�/7؊�W�Aad� #s�����4���Lr�gĩc6�M�xR~���*��P���\D���O�t����Š�lܥq`��� �xuL"�|�]����M���Q��J<ґ��;�+�Z[���eqW�LVg�re|��r tS�B���\�獘&�VmpI
��0)]wh�؆ݐ#��iب���VGD�����z���sKtSAz�\T�r!٣~�+޹7f�	��� F��w�Fh�t���q�y����d�t1���{�$!�40��"^6}
���i����5 �� �M)�H�������I{�9�"�ِg�&V�+�'k�`�&[*�,ݤ/�+��D���խN��2X��r�׈s����H�y���"66���ם�NDnԽ�îaZ���>��n��R�[8#91�G;e黈s�Ρ�"VF[#�� 5�EWo��M�2?�[�(Uq'����^��1 ��J��E/�cZ�'FH&3�W��r�,�vd%*M ������1^6�r���@é�f�0R_N�z�c��b�*'D���#��\�!��,�˭�(r�	5����"3��(�M���R��+�te� e����r��u��N7x�S�Sq]���ĘYh���Ӣ�Y���k�x�}�beςu�B�B59���0��
vs?�̤��D�s�閭��1`��W�)V`�G#�s����E�eVŤE����f�c��T^�'�W��aɒE̢�t[FF)*�X�1}kb��*d �dN<�n�Yf�b����ͦ�����f}%2#2�*	��b��Haɪ>`�� ;B�)��	�����@8�r�b���o��HjdoTT5����JD���+����s�0���p)-Ѹ.�\q�#������#��ד�Q(U�Q�]��D�+���k�ƯQ���U�$s;�!�	*�dO�j��z�J�M�X�k�ITq�2�bT�2#������p��h��^T�A5�k�g�j#��+���N"꧘_�F��L�B8�M���85�\=��� ��x�G3�+-�i���h�N��wj=�㙖�;.<��3�6�!�!�Q(�]��16�p�Q��W�f����<r��HOu�V�bQ�N+��&��y�E��S-�Cy�f�C"����M ���o��;%��:F�n{ű��d��
�1጑�b�U:��*I~��� �l 5.��ŭ���@��bҝ(�̺�mfVo�d����6`�O�_��52�k�v��ʾ�ϐsQ<�vO^��4pJrJf��Vu5���R3:^b鍟���HĘ��<#U�4x�ɉ.�z��� ?�^��M!lø��2���/$��k,����]���ww�p�P�������P�D�J�1R�R׭�P[��ŀU��0����� �� �����
���Zn0�Hr�$[�f�ψ�>�ph�N�8k� �Ă�|��h�Y��O�8r��~��}�����������	�c���Ҙq�>g��C��a�g�<*Ʉ/wΌ�� _��i� H�{`G�tK,�Y��w��~�Kn��}+7�T�Z����0h"u%\!3T�$ ���7��l�4w0�^ ��V�7� ؿ!6�g�&Vf�xe�"$�����g��s�s��{�͟'_#�S�{js8@8����A_�Z]��^k]�}���^W< �fx��3c��b�Uyd�u��U��F{)Q)��o�4���N�8�N��3m���pj��z����Ξ9&_��) 0eO[c�鶯lO�8n�$0����18��7���s������R�Ѡ�^�#3Q
�
�4�鵜��K�H�����4�d�b�(�|�IM hh���a�T�(p�Ms4WL�8	(?�9s��T�ƥ���0,�s]R�#t
3qٺw�n��~�9�y��m[5���
CE-9ݘ�Zʣ���q���۾}��p��?��׽�5�|��-Y��_���h�\���6��� r]U��^ř_�/X��'��_��?��������t�#�H��f(|��}��vRd=����"�z��>�5o��׿�?�3�x������6#�l��[Ġ�	4�($��^��gN�&`�������{˛���j� � 揃�rAV�[�4��C<��:�CA0L$����g������%r����o�I8����,�*2��/�睐�i�%�ϛ�c�v(��w���o��~��9��;�߿��	���#��u�2k޼p�оC��>��������K�����O�{Æǈ"N��{g�w�{�5{@9"4�s�K�Υ���&�s���qw�u������߶z��];���T=�IJ3;�x��&AŝH�h��Lڹ��[���o��7�����ƁT��� ��$謏��FGb�*�[k����u��x�?����0�o�p8�O�����8�λ_3͉HS�f�S�̼ܷp��h�n��_��^�
>���O���B%�t�u�譈~�_��8�~�z�I@�#���z�?�����Wmݶ���wV�om��C������ܜk�ns_0�B��p~�x�_:���S'_����?�p���{��y�,]��o?w�:�7҉�<D\9ڻg(0���@�E`��E[+W�|��_��?�-[���e/{�@_��x�⹋��ԏ�^�e��d�a�a��x{��wRDHz�k���<�����_<��g:6⦛o^�h���6lب2�3��^��h�ٳW�Cw5� �<b�y��{
�[��ˑS?��?�|�˿��G{�.���V�X&������S��Lx��R�ܱ����w�����'�<r�-�,[�z۶�>�XoQ����6w���6�%�/Arp�7��k�+��""�-V/��{�3��?=sMt��x�������h~C�Y^�z�<�fQ[���&�h��E
۹_A݇�>Ι3������{���۟y۪����6l߾���	UI�れ&�@L�X��ٛ�㒏KN�� /��˖-���o���'��w�7�}�k?���lݺ]�Ł��R�m�6-jG_IC�>���������Ͻ�oz���M7��߽b��==r�� +@�X�D+��c�;,�\2�=G��5���/��{���
1y���ov	V��aCjt��8��_@�?~x箭+W-{��|�׮\�~vA�K����o��ęӧ�ڵs�����{д�_���<�֢�|<}��1���ݸa�ܹ3�ϟ�������P����a��/��<>q��� ��|�r
 c
`�[T֜ ��T��W�ⵯ}�#��;�q<J�������O~�l�O���
�v�M7����d ���k׮� Eo D�m۶��-oyӛ�ω����xb��^ww��]�W�l���f<��X؋h!f��188u��E$�?{G�s�㈤�ׯy�������8]O%�;�����s�}�C�}�GFc�t�2|�幆\B�n��W^�
=�91o�Bز�I��O��?�����;0o��CO������w��w��/>威�n�u�����2�On�������Ak���w�[O��x.�����t���{���?g�l������+V��o���\xu���N/_�b��~/�Ϝ1ߋm�
�v�-
�?�2κ�X���7��/���'8��G�.Z����g��n�����1q]����_�)?wɌD�0�o~L~�7�ݻw��]�)���_�7����3���ǯ�~�����_��w��V�#�x���`*0!&��Dr��TAxl�}��?����W�?p�3��ۙ3w�l�'���5����5V�"�-��E�z�9�aO�����w��]��Ӥ�Aą$yk�!Ђ�L�E�z������O��%�Λ��}_X�t��eK��ظ�ɅC�N�<�v���`���թ�Km�XZ���[���ݽ�ѴNC������ �����~i�_|�����?��7Î����03���}����/^L���hj́k�\s͊��vow"�|��������{�5v&̘��M-e<BnE�RX�G5sˤ:�֯��U��������<������}���!\O�<s�LT�(��Q�eI}��|4�g�@���u����׮��Ng8�sϮ�>w�#����/�`�ɣ3��-��15�%!��~^ln�ps��m[��{^�WἸ�q��s��?��'>����)[6oz��G/Y��-�T<FRDӞ?S"*�[6"OOBDO:����o���k�?�����߿�#���w�l��P:u�Ķm;���c�:���V�<��K���Tx��O���_�SK/�;g��#�1�ʜ��>��?���+W�:�/�9����j��r*Q"j�y�۽k��ʁ�{gϚ�}�[����K��3�r��)���~�ӟFOj�"�u��3cS�*
x�6GhU�/G�t[��Ys�g>��.�O�����㍷^f,�����x�k�JC�'f�4t���?4o�S'MY�x�?��_����/>��10#�T��m޼�{;i�ܪ�vv����.Y�(A����~�G~�_8o�|����}���޵m����Yǎ�d�Qr�r�*/��ڪ�4q��ڪ�fϚ�sǶ���������,���#�ߟ�����}�!KLM�1�c� ٷg/¯�<̊�d`ݺu`*#�Z��X�|�5+���{��?����k����u�֣C��Vx�bz��RN�9y
M��\�L{��N�y|��E�����x�5���C��k�����֭�P�'9R$����\��vΙ3{ǎ]��4�Y�:b��-��GV\�ʹ�\���?��w��_=��e ��#�"3�}�}k�#����/}��©S&��a^�vͪEgk�7~�7�=���^P.,�I�4�.���?���9�8P2�N���Ǐ�%�1[A�!�;��:���k�X�>�����k�������0
.���rX� 	t��=b�qaE=�L���l)Ԗ�D���>�D)�#-_������y�����̕��-۴��}���y�.	bFm�e�I4�[aAky���@s�yϻ���U&C�~���c���;c��� �5GMc��{8�C^i*�l�ZdJ䊌����6mx��gϙ���~��Z�M�0���&�Xm��G8��&�����M�x-j�7[�ivY�����~�7�+��r��^����˗/��h]Bh��7N�ܹ}_��{��f9(�Y��/o����o��=�~��$�'L�7w�W	���,��X[%?*J��,Y���{v�b*����?H��d��O���#\�O$K|��c��͘9�R��GMԄ0���%Ke�5�S{�����ﭷ��������Wp?7�[6o]�x	}k<\�g�^�AdD�������$���ov�1#N_����g����<a���%̆��v��)S�=�I %N:ح=�r����ڇ*�F9PП��_�W���gϾg<�Y\X��R��bNA�t?�<��{�ݵke�j�*���رա@7����?w�~�_�[g[���^K+&�/��φ�O�aIp�n���p{�b�r:�VbF�r�X�F����&s
�_��_o��d��IT�T�G*�ΞdG��C�����K	ӗ�}�}޴�X���S���?���K��~�]�z���^�*L=qrŊk,F̢��2�;T�o����=UY�p!&!x�,��s� uF��6>�3��;���c��<u�1S�)rB��n5aP��w][RB1y����E��?l;�6[�С���9�u�g1�8H�J�ѵ�;�Ԡ >��r0�Xn<�
[-�a�������t��[��̝����<��rو���e�U���96���0�6Pm�:F��ɳ��8u���'����o޴��p�H�5�S���V��d`�J�s�V��Ry�$,N�<>o�¿��֭�,�	1> :�k�־�ANk=�<�18���e���4�a�c�z�Ey�f̈%4�����L��,�U�w~h�xlߗA&6j���w�Bܒ_�.���;g��ߖ.Y�c��?��O~�o��6݃*i����wH��<#:s����zZϮ���s���/2�Hh�]#����a<�i�c�o�.>ºn���o�~�0y
��&�@2�ۋ��wt����w>�����F��)�G�����>v�0��'���;����3m�ǉ{��1s~�Sl���R>**r�����8d?~��m���أN���CagM�<����]kj?C���b��ۡg�<#���.EfNج�9A	��{������=��g͙�Kȃ6�&L���n������|Y�W�hB�\|��G�ʓ,m[��g�9O�bÇ>���;v��N8�D�IE����D<>���'R[~a�JiC����>��Y���|�cv��w��O�;u��A5g�<q*��t�x�5������'��<q�'����s>>?m�>�-y�`�G|�奘l�N��-�4�& ��3�O{q瞌E�����}3�M�:i�4�����2�ǧH�X�
�o\cT3��r� π鐮��M�=c��3秜�s�����N����Gp^ʑ}���ʙ³cD&c��O�]?*[&c�&�}���VL�D\�6u��)�޴�V��!�>���|�o@a#���`���S&��9yb��)��zgj��w��g>���z&O{�c��'���''M��:	c]`3R��'Mq��ۤ�S��s��q[�s�.qV��)�'M8r����~�!Ƹ��O���&�<�>�]��!v��P�2�����;n)�0�o¤AǸ9z��iĎ[ �GO����y��)���9T1��!c:H�*(�c���:�SN�k�Kp���#ǎ�<u�)~?��J	��Ԍb���M���y��$^D��Yx~b��O��V�$����3�3f��_�A�*v�c�����zt����COo�1,5aҴ��>���{n��3���8��n�!��J�Tj"�&g�q?l.����u������q�k��J=�&�ޛ����]�efV�E���!�U��6�/�t�ܞ��V�t��W��X� �Q̟D�Y�VF|ipcݩ���8�u2��ŷΊ�3A�B� Y'�*��rT:P%r���K%Z�t�0#b���1�ԭ�uC҉��l�@��ݨdfR;��^ ����W�`r�.a�`1����}���l���%������$'�3\�+�!e�It-�D�.W@6ik�+�`���&�I[1��n�.��_K�x�i B@������j1 I�D��k� �/���?�PbĻH� ��x��S�5�*�$ؐ&iRg�*0��%9"`��O���Q��X�AIL-����`yN�;  @ IDATFFM�ՅT�d�D�+�}���ShT�b7S���b����P�?5��%.���s�g��E.U�&��a}�|���H��\�U�IBs�*��K �UF�w�������_LQ���0C<��[+������ w%zc��\�n�x^���y:�@�bW��k3]�)ڤ��**_�)1&�LM����|�	����I넺����3�L�Xھ1����Y+�v��); �����E�ݵ�쎇�QE��=��S��k���f�o5:�gX�J�3�$��i��.���Zɸ�ٮ���Un�S1��⍝�&��3�.;7���^,nmN��c����~��o,�|=�S��V�y�͌��>xRj���O���CǼՄ(�!�~�;n��t��U����:+U�<6�kg�t$L����{Y��S��Q㒸�x%:]�[�bm/:w��io=��P���l�l� e�O�p�Q�'6p�§r�{���#[���q�d2����[���鉋v��d�za�f*j�᫊�����(�*�;nδ4���`���̺�)/�R��*\��e�f-��1a�cvq��Z�\Θ��2/F�rb����|�:���v ��#�@��g���z�Ʌ�Y<.���'����0��������%��hE�X��l	2�ѫ��lgI{$�;,�%0�J1$r7��va۬E;B~��G�)P���FT��QŞ�2{�P�B�O	�)�'ՅLt��f�L9ps�.�n�na.�F�wt��1}���3�B
a�T$����p��[5��g���|�m}�7�>�}a�V�wX�Q0�����Wv���옘G��T��_���6�0���w���a趥U�����S�p0tJqJ�®3�&��S��T�:�-p��e��En~���7"Jl���ߌ�S-�Iw��:����n�t�>[�[�vQZ\�U sZ�E���F�%���/�Efbo{!.ɴ�4�Ж�����N���W�f�g�H�=�5N���.�n ��)����b���.ے_u��� $O����Y��1f'b0��1I�d�9��6��FZ�
>2�����t��+h�]��t$��:!^L4���ȋ�DT�x�d"d�� �p�Q�
d+�_m\����A��E�1�d�w_~2Gۇ��a��6o|mc� vn���ө�U����R+��W��U	�,� �V�J>�+�d���ݯ�n~M�i�m[u9�\t��*ם������*&�œ��mo2�-�8�-��	͗���㫈�W�ӗ�l[8{r��U�e�K�eӗm���˖�ƺY�k�+��mN��� 69(��œ����4O�B��X�_�T���W��Q���%�2>��F�RF�ĶY�u-תE(�����W���ec/��	u8��*D!�f/�����q+�)��ޏ���U� ����Mc�j�.!D#j�4y	8��� p� E'��}�����l$�A��~գ���$�W�'�������-�m��h=�=p>\��s!�4� �DC��NҶG�,qީ�p�����+��I��$�rw-���F���&��5LM"*gS	��0Fź~.+�� ������rt#��F���	gϟ�q�o�Ȋ��/��c�q�;�WN|�=|t����ja�t�ߝV�>�uU�b8Z�����g��9v��Ӎ�tWA��U�N1��)���[&ե�ͩ�X�?kp�ɣ'=���uZ���B��"��8ߪ���mϠ����7��/R%\Z#I�����0��23a�i==\�M���d�;8�����$!	>Hl�9ّ��a���w�&F�X�uƫ������GO��w�Ƀ}�O�����='��x2?󧞂�R:.��V�u��@W��r{&N�0n��%=^�n��7�����Y�;����l4�	����
�VB3ˣ�N�����~�D���qߴ��r���3���s�"�4�ȑ�ϝ���ہ�/ҝ8v�'���}w�Եo�N��c��L�|�ȱI��-kY�l|��rj0,bJ�M!������w�ֲ���`�;P(&�&�=yv��	�S'\�<��k �h�l2�]��g��r5�ͧY���a�xb�����@oߩ�B	�ϗs�c��M�1��B]��������Oç����8�=Sz��sgx9�x`�n^>uǈM�ȿD��n���Q�6�?Ɂ"�3��"��fq2q�fn ��̉���1<,�?�Ɨt袘i�|b�;@\�h�ߥ�o�	��+��i}On�<��ݹs֯{|�74������|���}Έ}8a���|O��q�wǾ��8v\"���q���Lx�ɺ�F4!��h�2�3�LZ\�^�������D��y<�������#���~$�rT�R��
H?�lor���7{�l�O
GX|0��g1c�v����7pb�"�+�bЊ!#$b��2��Ђ��Ws��ѭ�;vΞ53��
GF�w�4��i��|�r�J�+�>΍|�z��^�����%�@!A��,�t>�@�9��w�xp�F�y��t�!�'�*��V±Kc3��O���a!��q�樗z�BﴩΤ���Ώ'?�9������Ս8�龄O7���/6���Q'�<v�~�:80��aO�ʎ�en�i��0���{��`�ф���iZD��.y����z�7�4�bi���~O��!u�d�x�e�3��J���744χ����쁃{i�K�;��4�(��\��K1���[l`gϜ����3gL?>1��QH۶n��,�� ?zp�1ƟK->v䠊���@�Pr��n��4�=s���zx���G��d9��%s!7�EQ�^�	x��U]&�Յ�Deі���G�p~���ٳg�ر���#�a�cǏrJ��{HMb]�)gS'�0KD�	��9&M
�%�8���k�s��e릕+V�?���v{�P��0U�����_1��ʡ�'���� SǴ�q���ԓ��'^�2qױ#��͝=�o>^H.ĀBB��-�Y�[��`YOx�0��9~��njM���9�x3�9z�o�#�kB���X����b��E���3a⡃�-]�m�Q� i1z��)=��FO�#(��~��)}�(��2��`6�������s�G��8|���c����>��ᣆ�˨���U������5|PM"�y�\n���Y�g�ż�N86���e˗�ڵ�O���`�Y��hTDO8�8yɲ�!���^�I�m�i�i��>�:�M���e�\4�\��B0��T�ɀ��#Gqb��)�`�oڼ��eKBX�͂�b]���nႃ�c'j��<~���-]�{��ŋ�~���޽��uU���4z�{$�fF��,ɒlK����)?���$�PbҔginn|�ې�M�N�M�G��BnJ�z�/�R;��6�%K�[#i�y�G3#���������F����:���>����k���ڏ�V_#fu��}�}�ߡ��`�^��!k�_7ɦ޺��h�ԔK�6����<*H��2S�a?`!�B���4EӤ�9S�!N���pj����u��1��������67�d?2)c�d[Ga|��g����a�{�^ぃ�5�� 2�� �O>�bU�e�.�D�eJ�dDjv�~Pc��SU����-��ɒE<-:����kII3�<r�c�D��o�v��uWz�T�Ag6�?(���R��xn�}�'zzY'�3�W�G�G�SX٨fx�K� B.�T���<�i�&DX�޺����۵h~�]Q}�����"�C�.zc��Z!�da�+����x��e�
_�0u�A#����K��Y_j�6�c��V1W/�P����03�X����v��C�W����SӋP��-k�Q� 9��A1UNW)�x�B����SU���<+��F@W��4�����`5\��wd-~�^i�0���CQ^����@oO��Z��">8ןr��W9ΘX��J�#Zuu�u#ÃX��ojmO��5����NMN456(.HB3�L�4F��Kx�Xtn������ZWW�ʖ���8}B`)�R��Nzƞ`9��"	`lr ={_>(��1���Pk����N6�W�j��b��Xr����SA"�D��'v��udydt��}5�&M1��I\kj�#}W�Kݿ�4+���1�3����3����}�ǏZRun�.iz|eS�@�@��)�+W���U�	�`GϜ��:�+kl\��g��gr�Q0���:������E�mu�˿�̮�˘^�������&�:E�3@C�4�M~�,���%�z@���sR/T[�5�>�8�RS�^�Q��4V�R��n�0nH�X��EU��):�X{[x֠��fߟ���d��~ٲR�GLxpYL�%��*���Y��ѣ���ICȱ���6�dpF>�:���O�N����6��m3���{�joo;tx}C-p�M=P�*s����T�����c�1I��>M����w���7�|�ѵ��i�D�ƛ3\@(n����'�wu�mmk���w��nݺ��甉%ˉ�j�
�zN��f 9@R��U���:Ǿ�x�M?��}�[ooiY���x��1�ůDsX))�#��Ҕ!MTϒ�;��}���n�ap)����.�܉δ��聣թ&8�,�??K&��g����~����>vd��M�ٲ5ʥ��Ys(ݣ��q)�A�1��=�H��u�6����x�N�C=.]�����mF d2�{&�{9�g��������~�G�ݶ������G�\���r1���']��S��m�u���w�t�M+�٥��ú�������)@`�m�b�7�5����w���C�yӛo���RqC(�a*����t�
�3W��6*	DKl�b���o���ڭ���36>�.��R���
�������C���?�S1��*��������7$�qǭ71����NC-iw�K�	�a*�#Q�+1L���@ou$���{{������|�������{��ƟǷ�M)oii5������F0��sc ��~���Ma5��9E���������4N�~��Ou���G9� nhﴈU�+��Jf��
��۰ɸ�0�v�iL'�ӿJ8����_{�u��S]�;::>l�%�te�Q��X���'��5�)f�ɼ@U�X\đ�����}��ڷ��Xg3v��%�zɂ�V��.� ���W#K���ܷ��LN�+'�LKk>��_��ޛ��oz��}�=�}�[lI�{�Z�*SG7l�p,O�)���%8��GY�!�577�s�]���w�y���r��,�3�K2��t]��z<#��[pT!��u��U���c؛1x������wܶm{�M7���'�����K�9�b*��y�V`��:���4��s��;�>t��t�c��^�c뭷��u�:p����@�x���4/���ҭ���T��"�ռ��9��V)���]���|��������ﾇM��~��5�q� $+�?�0��Ī!XU��d]M;*��I�h�m�5���/�{�]�51+6~��P)�VC�?�b,���%֕��.B���V��xJ{��L.X�n�-?����1s�=�MMt�k��V��<���{E8���`E�lj�;mܸ�C��x j�^�q��M�q㘺��Uzĺ:N(\�\F tϗ�֭[��,aL߼jM���Sw�}۩�}��b�mo���w��.�µ)�l��-�-�2L�U��Lg�y�۞��Ks�}�=����l�B������W_}�wb�Coذ���J�nٺU;q4",��w�
\�i��I��--�֬i��?��C�Kש���o}˛-���if\���7���m�u���[�na�����+.L�ε����o��7�ti��W�nݼ�y������˹�hj��;w���
\���p�-[@S�ƫ6��ja}C�}������Wmh�:���oع�mc�㺿�ֵ�k;4n���ĩj]j/�P�GD��/�4l۶�G~q۶m$aph
����5ҮS�a���H�l޼�8�P1��Lmt֛p�bZ
ΘK������7nle���ֶ��������[�n�t�����m�����`�X�2k��-�_ӧ�p]��?�+���V��K�ę���s��!��$n��ڡ����ɫ���R��u��jU��ϴ��;n�g�쟬[�FV����k��45մ�XxC4"�jD4VGĒ{� ¹L�4�������a�.~2�l��;еZ+-T���AΥ������� ܯG�$�~��P�F������ލW��馛v�~�U+_Ђ�,j�U��U�C�^�-L7�����;vl�]�{����7��u����25Y�����^�K &/����Dz�ܸ�q�����_�v��S�#�k��]�Ȯ��v�nw���1��QԦ�f5U���6}��DT�72R�e�&4������Һ�����5K.W��O�$��T/�������W65O�M�qŦM���L"B� ���o�������wk8,���0M��G<1��5��v����ŝw�i�EZ(�L����ѥKj��au}V�I�BUM�V��8,+(F�뮻1��Ζ�u�3g���o��ݧ5&��7&�JA
����w�;�'ԈJ�� $}
��ꪦɩ�DP��q���t󓻞є�K��⥋jj�3�0�{v��C�M��i�I�� �g&��͍�ھ};*Q=�`���[nٷ���Ukٱ�nH��ɑ�/�� ��JL6���N5�W��6mڼy��n���BO2��N�$���\������пi�Շ��8��Ѿ��Ѯ�}�O>��?��,'�DA�{�n�how%�#ִ/�G%�]QS��/��>�S�=:��}�����������j�XO����-��y�޽�xTV��J�={t
"��I�~���?���?�szt�O>�7?��/~ed��0���zk�#C�Ԙ��ǻ̵���qVr㼧�zJ�����ڵ������Wضm�ѣ������[��놇8(��@1{��MgP_�;���^�޴i=����i�ɦȎ���Ͼ�裏��o��֭\1��~�7�������g�%�ZHM��]�p���BD=F�MM��if���1��ΌY���������~꓿Բze_�t_��������㖶�ɾ!ׁE ]�=���!|�����IP[W:����?|������ڷh��׾�'��+���w�֬�ypxh���5k[�=0]��F^a�i��H��:��o�����~��ho_5q�a�_�ҟ����_����$M�0H-�PD��̞<�F`�vz�x?��	o}ݢo|�ɯ|����W�?�5�0��*,� ׮]�BDϲN�DtA|qno�����D���^xa~�ӿ�ɷ�z]__�8��棿�۟ٿ��٢܃��`w�$"��ȋ��D��oع{��ᡱe�j���d�������/|��m����F�TA^�8 (��T����g��)��#Hil�MM�_�������/����Ͼ�и��$�N�rE�<��7��^�!lF9r4����&-D�������C_�_����vn����0}�m�©�g�\ ���^I���עœO>����|����<��'���/�?55b<��	c˖MZ�>����-���Q4�W� �<x��'�s��w?��~��������tyy.5�X���/|�dl��SCz��M�L��P;{©�B�?��'����������tw�bh#�,.aT�jva�QA(�u(�kk׶��Ԏ8 ��u#�~�[��f���/��/=�W�o�f{w��2�}��b����hx3's����l������2���4;���׏?>88�s����?�җ�㷿�K��;g9�[�ʘh��HC�B	pw��Og��ɯ�ZV��_��]O���d&��O��g?���L��Ƈ@`R���L�����@��Z���`�@�<b�\ ����?���;�{�{{~�w~��ǟXݼfݺ$?��Fњ��vxt�Y��!��c]�m�NVդX��nt���p�}����'GGͿV�&$I-�lݺu55�:��H�b9w��1���M'5�n��q���L���M[h���!lEK�j0H�Xs��Ȏfo��}��v=ݼ���K#u#uØ�ܻ���^�2\��Q��ڲf��Wa�k���#��/�1?�����MY����%'�h��[h�:`b����	X��*�;�����7=���O|�_�x��'_�����ʦ,��"�I�X�f#�)wFd�(⎾:| 8�+Z��=��w���}f�����Awd�Kː@ud��v"C�A��	|l��X�#��x�d����:v����O��:1��82��lpO��꯲���j=����[��g'��]��;�����<���ZO�К��C$$QOe�teJ���\����S&�aYmm[�{�����?�N~�_হ������oЂ m�x�ʨ��M�a���p~��J@zǆo����g>�oy@~����3�°�@�l1�r�����d����BU3ab�]����}�߬Y^��۳�ɧ�ä����ᑫ7o�4d�t��uYM�h(��)ǧ�����Ó���w�y�{���#{��k��~��8��Te�����~�*o^5 "�ohЛ9aRe��h��ښ����s��ר#�ԇ{��/0�5z�;��є�5u��e�������P�[ݝ{n��:_�t.,��=��x�:Gk�b9�6�8�����j�,.拦���Z�:��N̤����p3�Y#�Ҫ�}����1��I��;v�����l^&�(�S�N�8�R;40x�	Z�)��Y;)Q���2j��iC[��-'��q(l��{�x�.a���r����+�D�6d�Z����_'Ӿv���#�O�ԠI�E�$��hll��7^��[X9�]#y�I'c���qE��`ߔ�U�:�Y]m
y�g ��i,u{� ����}t�&6*�p��@_|���U�V5?�dĨ30L��ֱ��,\<�mkb*�+S5����@��,)��%ӽ=�˖�r|lu���u���,�鍑S�l���-m��|AXg�@Z�62R��B�d.�M�(s��:D��-4?��B�fq4�+�W�w�9<�U����W�vƎ�Ѿ^E�]_l���96j�uamM����}�w��>�{��~CU��Os[S��1[�fM�	��ɦe�J���p���]+��Y��!!�S"�V�o+Cu+W4��OF���(�(���e U1,-��]<Ԍ�v����m�h�̳cV՜�ݳ�y��fm����~���3�ҕ��$�p��Jɯ񙵵���������N���w��q����렻��9b�n�#�P5�ff4��Ub�+�=�t�z��gϞ�{���W�]��e[U�a�Ŏ����C�K�"�%t�=-�oY���L��k@�O�t�踊�Z���� C>�Y&`�G�������ŉ�/R�Y�`G���'k��ir��[ޑ��4�d�U��J�>�;Wh���G��V5E��ڵ��=l���E;�u����U+J畜�R�rg
�K{e�C[�]=K�V/����<y͵�ԁ���U-ã# ĕv���P�ԥO�R�.�X�a����Ti
�T��*���&|�to}݊ɩ���mr��.'DU�OEc�����8�d�F�/o�'$�GG���2�������/�g��"f�H��L����iv�/�<�)�*��r�ҋ*U�����'�Oh�zs����T8�Rqi)mO�R�\~!B3+��uMO��C�-�\�i�������ZR^��@(�:l���]	Ÿ�6BO��s�H#�nԲz�C��g&;V][�ޱ�`(>�p����߉��uR@ATY��=��B�fV�7B��n�n��fb���e��uZ�B�ܺ���̦� J���2cy% ����-��7�ֵz��ӽ�l:HODu�fDK�d�Gn�D��hi`�EJ:z��t�+g2�늳�`N��G�5U(F�dTP�Ļrݭ�\g�jjHi�Qc4��Eㄱ�|�������j6kK��`eP�=se����<ڸ�A��]�mW�v�?�=:>=6��	H8��b���t�s��p ���H�*P���+%� &�#5q�@�]����>K�1oI.����},碫�e�K�@Dӈ�I&�^��9K�� �̖�8��̲����U��3S�و��S� Y��|4"�Oo�ț�z{��aű�����(jO���^���U�DF��H���~�/��z+��$ǝ�6�z�;1/�lW�f����B�t@�4�|хIlms�*{�r�YӦ0��������'�É�;���@�w�L�mj'��C%�pD}Ҫ�2�o.Y���8�K\6l���c{�U�yh8����b�S�s��zQb���.T�F��H������(=Ǻ����ߍ,���^e�^�=4褵E�X�q!% �JI���C�n|,�.��r{յ�Z����	��E��gF�� ⋺e�	�ۂ��k?JU�K��(`�J"����qp&.��_�!ت����#�r���g˄�ャH�֭-m�'ݧ�j��gݨ RRw�	��*����G�{��_�1f�ʪW����H�c��4��.�B;0L��r87���E.pzi|C�j@V��S�W_��?[�E�1���q��a�R3���%j8��ºHHF3�.�}Oi;thddQU��D�@q�©s �m$��Ua�0���QT����.�pkǘX_[�F4�������j0d� �h)dA�|��+u�i⳰�Y���̙����X�ik[CK^���0عQ�bR&�%s�J֏�4Q�c�B�q����$}
2�U�%Ƒt��G�f���|��+6�њ�M/�oBI_�W�D&�^%�E�|661:���(i`�`�W��W�L��CqJ�j�|�h1 D�,דS�uV/�7�2��f>�[�lI�D�w@�>�˟J�׋��e��0�h�2þ�#�bIo�V;�˷��OE\V��V5��d_�ƙ��V��Y|��hgu��~d���������vm�C�����Od꠴V������5	q�Ӛ��wqd� ������C�C\�/��Ϥz��� ��W��-7�Z�������N�c��(��N|BG��`KO��ٺ��T��2M!8 ]�u��KQ�Z^���T��O������7}ݽݾU#'O-���/E�Ew���X$K�ǒ�3��#��Ъ�t���j��Ƙ>?a�'�n��b?�A�6���I/�R�D�<�S�-0r����¥�Ї���e�e{��߀&�H��%�|p�Q��Wu��f��,MNa!��q��xL��U��p͒��K�1�jי�<:HD��/J3�H�rUp\R
�#�d�R�:.�pr��_Ư|�P,B���K��x�� 2�~!,��� _Za׿Z�6DЄU7J�U�\y�қD��PF�2�!�%HJ�nbJ
P�A���$�#>A6�9:����,���42ł���9�2p)u�ϫ\bN�1���"��V/�}F����_�]T0]���4�o�`��	�v)���0�+�g�\D彲���g�3Jp�;�τG�҅4�H�0yc�-� ����?�`?�}�$H&T&P�J"{_V���:Lȫ�`Ѭ�&.�	[%���"�8�6�_��D�U\�$�JW9��*�� s��BE�W."g�+1eO�`��j�I�{�G1\�^]W�9V��.��|��v��(�c�kzu!�¦$��y�T{V���en���5��ǉ^�,���Dy�ΜNXDJCQ��g���B08Ϙ��������z\|/[�2o��z3-ѫ��3�yR/_3�(�F�P��ŗ���?��%��6H C�5ǉ�<:��%b�_]W���dL:�*��f�"��13������P X*]�1O�Kby����E��X��痳�˗���d�LZ�Ͳ\�7�t1-�9�⒕)�rV�Re�T�zP�y��D�M���K��+ﾟ(�]�S�kQ�̜S�"�2\D��f�y95���O�N4�~�D��)ܝ̐�r`��i��朱�l��I��xV��q�!3�ˉە�^�%V&��K[1�.5��3��JWZo_�e&�q��b�/L�c�� �"O���\���U�$�+�\G�	B,9_ᜋ�+��;�!MZiRK#s��y��>/5>7S��W@F �2�f�N�jC�������h�Tw��o#P�H�>��[�$#��E������QN�H�W"�c�I^ֿ}^3�e��6�\n2�sÉ�i�q@"�������iI�X�����jn�$u!�0Mm�rŖVz
�s��&s���#�[ZI�e	Ѭ�[:��7T&<�(j�$�4V
�Ǘ�+e̡@�����\4b��\Λ���JA��'Q�y,ǔz�$��YW�g:�,s"��^)��y8u'�>]�+CQ���e�X�E���_^����@��h�|i��ъ+�H������UBf�<� ���Ť��4-v&=V�RJ��Q�|f$B�̕�Q�$�����8�}�fY>�B[�d��,���W�/�Kn��@�L(_�hz=�����oV՝N���i꜎˖0�����@�{i�}Ũ�'3y&����ј��>L���y�_9��.�_1�_��(�/MQ&�J��H�w(�^�˼���ų��U����q%�a�q3�JR�J�'܈cư'����C&]y�,5Y2s'��_���^�����'�q�3���h�W�@�2r?"�w"�9f6v�J������	Ɍg��6Nq3���JeY�ʽ�{v;��O����rc���$�-_j�])@!���r�1��ޙ�BY6x��Fl���+�Ɨ~�����L�W	SY9��AO��W 7�o~�#��\RX�>aJ�/�ch�9�j��<��\�J�I���j�8�P���W����i�LS�g��cr�˿�,�!����1�<��Qi�w�B%���%���$MLr$�����|����\�rd����/��� ����.%b��"p����/6��03X�� �u��r��� L�R��'"����M xT�s�9Fͪ�D�ud
z��5rD�.�􁇌�����H������&}���K��;s^�*ق����S���!��Ǒ��X.����=6�~J�ɺM81>;�-�H�]bV����oaW@>�ZN���'�d>���d���+����ח{F���������]_2-��n���cCg�'V41{������Xg���wpd�����C31gC	�����u���O���ծh\�xQx�ɾQ}mc�T�d�g��)Ց]� ��C�˖,s�5*x6�����W�~�TD������g��/_h�J/_R7��ֻ5�Ν��g�v�⥓gk��O�M�V7@y��9�.[RÝ��ș�eub�P�M!�-���9?�H�D�%5�k�F�T- bz!*^�Ό�
��Lmj��5* ���X�%-X��Mn-}�j�\�ҫ�%�y_;L�2!�&�,�q(�z���ƥ���~֎�uc
����h2�sL�+w�ʴn1�u�_O3uv||pŊZl0��R��F�$�8)����Y�Z�kzl�W����?s�"��U�tl�1FT�s˖ħ�g&��=s�Ŀ� 6�!i�@�X��fT��aɄ�V	|�=���h��Ūqu�[}��������{�s��:����-JTW7�����2�]��{��vaί^���}:̂�b�o�-��da��.DoX��{��Y>��k�!0��ٲ�Y�����,�2Ss�ٷ��&3|d<e.\�x�����eK�kՉ1��P�-�p�8qh��k���!&	���$G�� �=k�`s$�/J�-3g����S��O��AG;���'������o=|� ۤ8������
Z����ĆŐ d�X�`2U��L���ifX����k�[�ֳ�Tӄ�t>wf��=ǥK���rA�����!WNLh~k�ZY�h<}�8Gc۶]��}� !p�1Z��I�|N� �'z�FP��A@A��u"�3�e�U۶m8=4Գ���O^^I�O�Ѹ�>sף0�}a�\xN��9ec	UfG����kښ	�@���gq��jcZ���� i\5Mff��yG_��z�)s#j/"�ڲ�E��75r��������f"rhnؒ���0�1�P�9�@`�+s��AV}��
��ܜ�m޼�y}�0|}�+�
�GGF�I�j�&�y	�ŨHd�S*#ʓS�ͫWLL�9��w�iE�;�[��t��^�~|��ھ�}}=�5p@��G����G��GAc�Rz'Ό@;<��O��T���Յ��,���DrA����DsssتK�'�A���M�_���������NIb��.c1�1{�L������G�x������cdhptd�Ecl��w����M7���#�p�;���alt�ر#��g����ѭ���C_/����~`{Y��� ���� ��{���胷�vc]mӑÇea�B��n8~�U��c�*-f:^���kf]��?|� ��<�����>������޹c�vΝ�{�{�������);��::ڎu�c$�����w0S��7nX�E��Y�6����Ho�u�Z��G��O>x�C��y~t�=�)&ukY�ck+w�ӽ�܄��.�E��镫�7ll?q�Hht�a����1�Sʏ���ʯ��Ν7>�BW�1�A�������~WqW���=�dq2�\�p��Y���������wl��G?����S�L�~�;���*��Bs^����&�[�0�r�U�h�DX��+k#����XyםU?~���護������=o{㩮�cǎ�<�	`B�%�k��H&7���aI����pv��2�"+��"�@{�i���k����w�����ٸq�~���c�త̭�t�
���澾���~�b;ai�uk��։$��X�?�����y�?�ȇ~�Gnݴi�={�z��a���	�ܣeLQ2'�����&�a�H-fÆ�'�N��9,�������{������|������aJ=�^2,���5�Q�UJ�����'V�n��u���ԉ��na��=cƼ�o��w�֧��]����GTF1~j������,y��-�-���t�>	���\t6����������t�T�����ah���g�Q���M&?&;;��X}�Ɲ�{���u���ӣ3Yv���������UM,(���m�c�=�О��h?�?87��O��;�C�N�&�p$��{��Q7:2�_߱������?�6�I���;︓<?��S�S�Jr.�]=z�`�G"�����8s�����8���=���p����o��w~��֯k�:�uۭohiY�j'O o�ON��Y��Nl�x��	��{�ݐ�{��xd�k�~	���>�����?�frOO�C?��m۷��::ʈ�h�W�#�箓Ǒ�`�c
��bx���g�G�����+۷oy���������otڶ�Z����{���=��?<E�8�i�Y�3��0>���<� 9��3��c��x�}���P"v�]oܶm��~���Sȫ�N�3���5��>)�!'OtjGc�&6B��~�O>�����_�e�u۶1�o�ޣG��k`���4���G��ccCz�Ĵc�Bb�Ow��H?��z��;?��O�a�/tnټ鮻�<x��������՟2����c4�ę��	�r}?ز���W�����cCC}�l�������|p�ڦ�ӌ���Xk4��2��,�ED���|�אRZ�ގ �f)H&�(mm��Q�Y���^�g_���z�<�|#0+lh&�bXR���t`F����z/�kn���&EY�T�R�c���'�$N�^c.n�dTg%5h7�Y��+�<�ʳZ �����i��uBb���{�i��`"��	;7���r�>�$|�aD�>�\A�?����(���i���o�m[��X�#Ϭ_��������{��u��>yQܖ-[:�PU���]}��i��?��48�P���#Gr��w�8�Ei�+��)�ڵ�d��D��  ~IDATso`��������=��W��y7mڤ;��j�Wug�����BH�Be�S�ݻ�۳{��!�����F�.�R�%�Ǆ�@wAw��Xw��v���FQ�.Wo�����_��ߘD�B���r�VPD� iF8C�����y��nh_�F�����/$.�f�/��/�.��fGQ��95=�B;t�`�i�1-~�^x�n5�;�J���[�n�`h����!�ѱ���z橧�esp��մl�1�ʱ%&Wo�B�)��<y�UITBE\p�鳫�Z���+a��ׯ_�Q�Iѯ�묀r��E �P��K��Lt�z4�nni?v����uU��a����S��p�E��t�:�F����kh"�'CD����BD�HN�һ�b��[6_��?JPy��?׏��e�̊d�����������E"�;�4��P���d�;;�c?6T5��%KFޣ�_WG��w0�#�(���@@Y,���42�/�Y�v-�[R�W�V�%�2�S��A�t�&�iE�����+X�5�ĥ�����X�V�"��c��0�0X	�PM������4+�,s�j��Ŧ������mPA����M�͈�;����7S�����;��:�#s�S�B.�	��n��'AlCZ�F����LCw%��T������c3�P�c41�Er����"O��Y GUA)��ʐ��oM�e�,�G/��Z��{E�c�0�yaJY�L��Ġ��B�X�L��1�\J��h��ϴ���'��}��:nl`�:�Z����~,x ���F�/[�KA����A1E?�m<C��"L�V-b�rt�ɵ�t��0��gR�dj��%Ń�{!�f ��g0G����}����7'O_Ѵ���3�F�IDu]%���(�IFE�(��(ä&�:3S�da�l�:�g㋪X��U�gd��Pʣ�~Z��l������kM����fY�)�҇џ�Z=1=J)� �1Z���w�(��ҵ�r���<���f��qswb���N���Ъ��O�0�-��w�:w�8U>�Y�H �8�d�JFm���#L�+�ȌUՃCCe�o�Db�׳��Wg�ϳ��S�n��FW-��n��y�,&���L3��)���r!ɷ��]1D���N:ǞK���y��ޡH�*��D���44��D@Ʌz���G�D�_��B�5�h:����ںژ|�x��ˇ>zozA8��o�v*���� >�vO��B�B��A��c7{��f���LH�k2���Od'.���.`�) &�a[ZV�YiV��{�C� ?�[��h)��[��
_�#��k	`6\�tE.LKś:#&~�t���ڽ�O��C�� ������p~��R�1���Ī�-�0X�]����;Ģ���R-�pc��ׯ�M���RѪx����<�h,�_�XbRR��u�YL�6K���� m��Ǧ�W^��V�x�giLf��@ưcb`��`��f��aƛ�d%d�A0�*BXYI��j3��drz���Z�2����:y���Ne�	Ln-����+@`H�b:�g����x�cW�>�k��;��Pg~ݧ�֊&6�'��[��[k�`yI��i��f�U�)��E���aM��La�a��B*�>��G% � �؆Oޱ�&y�^� ř��`Zl�Qvq���'/ށc��ر4mU��TxPU�/���M6e�:��,��vs$�v��j_�ne�����M+���qH";�U�W6�Zv����i�h�d��ݼFq���~���Q��}�7*���[��+'xI+�Zc�ɉc8�<��ϣ�t�~�0�\��ܘRc`�C�c��:^���+&qӖ��S��*��*a�n�hi3�+�	�K�����2G�����PAr�}�Dǐ�N��N80&as)h=��Fs�v-��GҎ#�r��������/mٲ����p��L��
��cqin�s@(=�/~�\��b�T犌 g��RJc�P��E�)}B�"a0ŕ���"P�o�`��┋�2qRx�vE�����O����V��e_+�+ߋ�s"s�[}F�j/�H 5�p�$��ť��H�?�^�2%T�Ϭ�*�Z��w����f�&T���m�8QLʞ���LE}+k]�`/R��h�l��"�m^&f�Q�Ee&�"�4@���8p ��5X'MҾV��Ȑ��-�rh9\	�bᠸ+D�|��^�� �u��(���s�9��̿�[(�U 1ߜ},�
�*Q��p1l��" W
�K�����/������R�j�ꅠ��l�}m/����;?Ή�H>/ʳ"A�����3�"�*3�1��|���s�/A#s`X�<�oL,�0*sei-�Ae�<e�NQ�%�w1��H$�:���\6�-�.Л�^Y�J��c���<��U-*\@.KQȏ�[���[����m���2�xz�"�= _ɲEA34)�R ���os)s��%�8��o�,]<s����ŉ��k{�*T`8+x�t��m��"0s`���Yg�.�,k=̙	�F�1����-��%��7iu����bP%���9�.##!!f��D�b�0G�R���X�X(*��X��`���R������U����9GQ�켗\F�o �r�����"/QD+�{1�
���rPzr��.p��_�7(�%�����].�Cq��Cc��%5���f�+�.�r=gEW��bb��$�I���h8��rRB�bi�vЌ.�%��+�2؊���7����s^]�Q4���E��*�PD�����K@��P�3�9��f���,�O]x��2ټaV�,�,`f��MsAd��/� y�{G\ ���#�E+�'(�JL1	���&K�]�f�ĒU��Y��x���n.J���(j)��oo/�|���B|��N͂@x�N�^��襹�[K��H�[����"�L_n�"��bQDz=��JP�U�x���/� &]�wn݌I�-�Q%|JI����� �.R��}VAy�TưHs�@�z�A�3�k��5�\��v��E `�_?��G�ǽ��$3r�~/�j@�`&�XB.��fs��ސ#1|1��p;�'O�pV&����8��K흛=W;�4/��G���q���`�|�l�-�d��9
SQ�y��DʒE�TDN�.�E�p.k�%C6p�^ )��)�2q.�H��0���D��2���sY*��(��qv�y�DE{�X	A�
�����9Њ���Z%�$���q&g�3/��yVU;?�V[b�O����N<�E�(6�|@�)&=�Ǚ�H�9��1n��n�2X�V�l���L�؆����U9f_�m3��E�Bg�GD�����ь�������" �ΣP����i�r��A�?n~*(���|�j�K�͘��KE��(1J�pJ�<�J+��{�E��k�p��%t�%z)"�苣]���Qɫs�%q%�K�M�f�G>�-�(�����anМۈeJ�sf��}�ץ冔:�B�up$龖��X4q�fn� ���+�6���O0̺����1�h�SE����x{����}�r���*�]<�!́S$� `)a�s��K�_�)�,��*���凁��^�`�)�cZl�|���g'/P���k�/�ʩ3�E�"0/�K���b�s^hs#/�S\,���<ӌU]�i.�%T!���U��_����>]:��������C��[�W������& /?��{-Y>�1u�gwQ��}��2w��+xMR��Hb�s��*���$e�T�
^a
�9�g�E�yB3vd5_�0�W��B����*���<�Ɓ]�oWcR�c�������
^I
άҺ�@,�
�'5r
N1Š�J�{��+x�Q��Qi���4OXd_����d`�ly
*抈��x�Ju_ ���|Ro\�?Ikz�V���    IEND�B`�PK   ��W�iҶ� t� /   images/eea2c8d7-d880-4d78-8cc7-667d8a2c86d8.png��X_�=������������;��-8�[pww	�����������g�V�:��V_�Ѫ�2�```�r�����``�p��>9�?����8X����:rVJJ`l80p0ȿ(`����������f��i���6��7?����_�Z.��Z��``�p( ; ��68$X�?q6  ��Y�!��w>�?mڿ�[���i�����``(���SQ�ę���q�QR�7w��bj�df�����>	z��1?[���y}vpt���������JA�7������*����%7�@!�@FF&�baů.)���'!
77 ?+���'�'���5++������������ԋ�ѕ��A�G������f��H�׳������?8�������ߙ]�Q֟Y�򰲱 X�'�����"���w��u��prpr� ��[
ssqqp	��'��
U[/KI�ϖ���� �!�O�*��ܴ,]���k^�C�_��1����L�O&�`�j����l������}'��N���n�N�V���.�n����Aհt���?��l�����7�����?����w��w�_C�U'��|�W�turp���������O��Tm�ܜ�,.[s9G7K�˟������3�3�_=u�t����C�_��䫸��)��������u�]�0;������������O����R��U�}<������;�0� �v+a�{^yg00Q09I1M/�·f�E����O�|�?�w-Ɛ�eU�R�Q�5�H{�!5}Q��4��/�:՝4�� ���6�ov:$����,��M ͳE� 8=[p2��r���$�ժ�DdLb����Q#r����JO����е*��72� z�ǻe���H��k��	�(����:<�=y"e{����&�����=��Rsp���%�4�$\i�Ꜵ�ʒ�	w�޷/���d�\����{9�{n�㋒H�:��_]��.��z�U���"fK��lo���&[)#��Jg+L�:�i�gA�6N� '�O�ݘ̾���o��E��Y�m���79y=2���{�����/0��g�w� ]��q��%��UA���eaSp���:+l��ޡ��H��+{�3�ZǓE�>�XW���s�g�k��˕��6|hHH��'8�G+OE�L��1j�V�hђJ ']�wŎˬ>�Ng~0���V/"Ҽ���H��̳W�paXgҵ�
ʒ�@z�q�E�����,<k@ �e������`� ݺ�������=�	I�M�ƨ6���)`�W_:�WٕNǼ㲈�ƳF�|òC��N���|�����rT��P�Qǵm��p�nTt��Kp"�k������Z1�kqS��?oW�����Ͻ]ְ������Yx�.��Ds���d�t�e��Ż;��Y�<i����ǆ��>2�t&N��mb�m�{o�<F�T;���\'���҈e}i������%�>��@o��xV	t�U���'.K�S��u2f�MS�3J��JQ����ܚ4{���c(x��Ŭm��D�������;�Ҥ�ц��pZk�^���v,+�}�@y���V/���',��v�����Y;�&B>��wO6�O�JO�l0�Q�.�dBI�����C%�ei�?3��u����,�G^�0�C�����W�m���F?�,>�D��pꏫ�rB�N�Ԟ]k���&/�|Y��m�?���y��d�0��~Y��ɗo��2"����|�c���G���@�r���i���R��7�����1e��or�������y�'$SF�n#���;36�!�hUu�U��wu�p��<?	�y7§�f*�y�<��H�Ջwϯ�i��8�-��I���/nP�i򸲡;����������hU��$��n��yg��[q�A}=�g��R��̕�6ݱ�ԥ1�s(�G�E6�B9#��9׃zc4�����Uǚ<:�z%��;}=dX�Yg[7^b���.��#6���KG���7� �!�s�6G{�+#��sCM��}*�<x{�w竷1r��S&�tW �$��E�۩�Y,ī������O�Ҹqf�tO�>,��p��[�}�SB���n�+
�F:
�EΜV�<��$��܌	�/�ϐ�lm�������TI�է�\	���nKYe�̃o�Jsc�><ӠL$Sw\�w�l8�-�
�IW{as�!�dx�v���5NX**��uU5�E#^ �^ �E������c^�m[�>A�����6v<8���|;G,�%!�{.K��xR���@{���l_�@�H�|m��;�hS�_1����R#A_=g�;
0߿V�Sj����ݗ��j�`�o�]�zu�ZR�Ą�9��a��s~>���SP9#�YPzhEڴ�jT�����f�@������Jx{W�O�6�֬X�5/������y�Tui:|*k�mݑ
k�Lg�J�n��4˟{_�(5j�~݃�$��@4�V�G���f|
�_D���j��@���8�	���K�A�����b���5��ݶ�B��*�T�tS��b��O��F����1��~��^�l��)��T������m��f��F|L�s��
��
4�5���|�DR�z��jD�6���SP3�����d���tF�g�.�/mv�vqh�7�t_���Ѯ;�f�{�ˠˉ�w��I�}�1�����~��~�[��O����1����q�=��._��^ U̞n����-���7&J�F�(�O�0~�����3�����.<�b�o�,͗�/>�R
���2k)u�����L��	?"�v��\�X*x�M5�LwM.`���5s�X\8�Q�T�]�D�t�ճ0�'�EXh����цK��V�r�D��,�]��cڊg�[�j
��	u���	��`#��r�D�fS�t�u�mWӝ>�=���PF���^���qn�C����Jԯv�_��j�`n�l��a[��84��kd���D����MiB�=��f���oC�^_)��2��N�Y?�x9H�.���Ҋ����5w��]�HҹT����yi��G����i.����̆(g���j|���kvجK�A{B;��z�<�9���#�QA�]�h�����䤭��2��>C;j�ڏ4�X���z��-�%q��k^�ʩ�f]�,���	���J�W��?��?���2MB�h�R���i`D>p�!��ݚmq�c�}�2��{�έ����Sw+˥����O*�����U�����0v�9Ic�҉����wޘz6�]p�L�ssؑ�L|��i±G�~��.$T�K�����&7f�m�b�g'���eU.WX>��;Q��?{��j~�BY`��q��K�������h����ڹ���G6�И���8t��$�-�.h��%|d3n�����68KMYcUs,��=1��z����}�Xe[�X	���D���C��$�����4�<��3��;Ͼ���}������=��tW�������I��UC�N�Q�5as3*s,o���4R���r� l⡤ρ�J���F߾EO�*g�(�0:���'3C4�U���̯&����b����tW���&z� 
�r���2Wzd��%�;gz�9%{i��Q���׫��E*���n>U]^|�z��}R�e"�.C?w��\c cD�'��FOJ<Jy2t$�Gq7c��$B�h�����;m��l�
���3��R�E�O�Z|��	����041��8D��eU�O�(�~��.Y�����l#O?_���zQnH�{(f�G-��-8�dwaL�~���5�o�\7������Xgh̫�Bq�j�	�\7Pp�y+�qt���s����}�wŘ�w�o���F��@o�;FI�����n�����0]y����*!=�4��-HY�jBP�p�_� �����-��,�a�ޠq �d�^�o��e�$E	�u"�ܡn)eI�h&)4�>��G�B���˔.��RG���EԎ��`s�o/3���L��8Ÿ-f{��a%��w�O�3˺	[�} �1��rNN�E�e 9F˺�1h��a��v�4��Ǥ�U����lZY�R �S��8�"�A����#��o��A�9/n �A������������ه՛R����n��h<��S���w�y5e�ј�b�T�n�'�Fn��8��t�n�#T�m��O`��-�"�m�+���E�S>i��$B<ѧ��u�B%��������`k�5�쩧����O��a�-�r�=��	t\�%x�\ך<r@��kח"1!���vO{y[�<ڿ��ې�����{%t� ���K�e٥qx�`AK˻�� R��q���E14[kk|#)P!=ö����z�i�")k�4�}��j�Mg��|j��ٞ�H�*�t�,=5<�0ٱ���6���ivd�ҋ�i��*$-z�i���׶�G.�1����2N�Rڛ`1ۀ�ˈ�����-�+����?�6������<��\�X�A�������4Z�OD�u��i�N�M�����md����M޹������t��ry9����P7�o���C.O����}�f�������H��lMջ5��Qhc�!BǪ�O�(�} �P(`@���[_��(�?A����R勨�<����_�g$+=�N8(~5��K�wSX�.��o_���H/�8�j�n��]k�^Vc�:��'ʵ͚�ݍ���Z/�:�h�qxＵJ�����b�,��P&�Q	b�=�=`�z^�����O	Tj�V�����nCT'�M���0j*e�H��^ ��(�40��怶I�(�ƪ��[���B�;g�{���'�A��)ke]�%+6}J��+�*��EFE�[y��!�m)�xS�!�	�d�_m�$��У,'�/�A������"x(�Zj�(ْ��vn�Q	}��;Ӽ� ����T�+j�H>�ӵ���ל̌C^R!G�&1��o�_�3�)n?.���gb�P�ApϚ��f�m�� o͞��@���&�����7b�	�P`���#Dl=~�����FkrT��M�j��k�BC'bv;*���^)�{��	@d�LtJ6��b!���:�
&���vnҼ�2�ʌ�c!��~M޸1uz����zQ�-6�G�:@�J->z�΀Md1��a�!�=�Ez
��7O'�^������A��h���ʷ�j�0�Lz?-�Qc���H9*EN��Z���!�@
c�әI���ϔ�L�<jUe#���z1\7�V����ex�q��Ħ���wa9�-�=B$#�"R8K`t�����/BN�!6	jqc�����z'j�FN|�W����ϔG��d I�F��l{�}b�~����0L���^�4�o��z�%�؟.������TI}*���Lpݐ��ĺ�*�Y"�|���T�p�H�M���� yCFx}.�'�hV�G�&C�[60��p�#(}e%+�ʡ%I���G��vs�Wc��2�h�"Hpg6ɴmC��5�=̓ôB�c[��ݍ�D�:۽��p8���J
뭺(��H�yE9u��=%/�������&dl�^D�Q�>�����ޚh�˛q��%H��K�T�c�W���cT!}� ����R��j:�b���bt+t[�=?����������NulyIl�ӐE����x�}�:����]1���2_��(_^��CТ4\�\������JĊ�����tt~�:;�s�������
��غ�>�2�W�\ߒ��%�]�f�d.ot׋8�G�eG�7s��4D8�p���3bZ���_��DHS�mRf��u3�pZ�1��q���z{��}qk4�?#!-�p���@�#�k&A��?<�b:���~�ِ�3-�:E�T�l�,b;��|��s�G3;H����E
��o,�R�:��C�,hjo������	�v�_X�_�Ho�)��E�c��>J�N;�r���"m�͋�$+�s�]�����@3��a�3����5?(G�2e��FcȐN(SV���ًyh��~��R���������3Hxu�y%��X0��aH��h�����f��rEXrVM�^��< qt�[:��v�34I������Q����ĭ�D����>]�-4�m�#^�M�>lP��[�
7���EM�k�L(_o���/� �Ʋ���j>��?�?tl��Z�J;$�����T(�oV�<g�K�U�\�_�b���B�Y�qU�n�"������8�b��N�_ŶkU.
ҏE�w��+K����L��!��A��h��WVI�6�`F��|�G��qݽ�+7��;�0���8����uO�% 4>��Q%��Ұ|o&l�9��)X,�G�L%�lmd���y�If����^.D{g)���볤�oaN���`�i�t��Pn}��6QMP
���b��v1|��[$�� &�4��i�im���s�A����Fߙ��4���fe��so/��`�L�'�qx���_UH�4��i*;�F���[p�35+C�К��༈֕/�2"���o����"|խ�����e�[��~��֐>63t�:}d�h�I`��!���lv��[a���F�������<���Ȓь�4(G��^���,Fz#瓚;�1@8�[�J�A�y�����q��C��1҅cm]�L��9&)R<�>{��2c���Eεu����E�q�!AM��ow��6w�|\���X�k��|Q�Vr�.a����{��yq�x]]D���'��ޅ�J`<2���z��ɏ�����/��UW^JJ����r���7p�ß��0b�D������n�	>��B�7?>YR��q�ښz���	�l�	z���b��g���T�PΏ�ތ�(Q<���ؽ�m��J��	7v�8 x:��L�uU�[Rp��@����	 ��J}n����gF�I�7W'%Nx|��4>j��m��pc��;5#3��UAHF3�WS�_�3V
Z�5���!F�[NF(���x����m��f��i�.��Ҏ{[��<��e0%)I-j������:�s\���j-Z>���wK8��;X1z1�+E3������� ��K��qShyE:��+w��U\�<��6�e9Yת�S��K�2!�7#�E�PW�0OHx������d��*_���J�$V($�����2yS/�ڻ�e�g�y̗9�b��9����h���5q��L��x�+��@-6A�廽Ox�
Q���gb���-�i���G��f�Z�[����#�`?e<�(�F��.ʜ�����?e�,D��q�-��*������aٱiҖB���v�͸���=A���G�mi���X�"��L'��Q�"�V�Ru[T��l�H>3Z{>����[���p�e ]��K���p��營1�5�Ƀʯ/���&VAIh�s���A�L�D�.�G���`c�����;3���V��{ǵU%;=�g̝'F{�M÷�C�h|sX��/��n�3)h��NI-{��k�$��ε�g+]��kGr�э�H��C���~ūG�-�e\^�3}�@p��ٚp?(�vΞ�\:�Z�rz�%��oC�������9T:}��꽣�-��?���å�����u��11q����U������E�fk3������L��5'����z|Au�}����F_�����Ab�4�DmDTJ�n��i�*��l���?[��x���hVD��>���ǂB�q�k�*�}�`�NlB�T��F:��kΈ�G���5�E��k�R����t���pqI�y�'�q���W���s����C���O��e`0���aCkB͒J����l��GM�Z����D��Ӈ�כg�s�վc9ˍs��In�>�������:�x��5�i�\�${z�DY���Cۜ�JW�U�A�#H��H\}ǈ�k6�E��l���7�c�r#AV��H�EMz����>���uKu��5�eBg/�U<�%F��Xm�������ᄥ�:^V��Pu4�?_�=p���Ҙ��1+�6���u4����S=��kTNX2Fgr��xYX*�&<���vt(��D`���%�B���H���&([�1���ӿ��^����p\�>S�����M(4v}�t}䤿/��/���#��B/Yb67hj�KC���ah�e�/_�A���4�I�!�麵��wv�ά	�܍��+�Iv��vݞ���|�|X|�	�[Թ��e��C	��Cn�Ķ�Jhf˭r���f���ko� �4�����5?aQ�3�X�{lKF$��d�/ʫ���3�����/zؼb�ϑY��8��!๲�yU�a<˸�NܑR��E��Z�q'��!J�� ��iU��2�g���q p�j���=�)��,]K�3�U����Mv��[�Xjװ?��N63V��
���)�<�жA���Ҕ�;R�ҟta�I��{�թz���3�\"�q��'P���L�&�%;wj�	�9�����&����+iBGخ]�$����v�	�Z�	2'y���0EWK�Ա6֟��?��|N��
|yo�x��|G��w����pR�S�����*�z�X9���#2�n8��[�-$&�8^����U� 2-�Y�ҧ��5yk�y��e��c/3�LS���pq�Wı��՛ه�������bQ㶛�<wR�!�w���͗����@_w������&T�.`j���,;�ָ|iߴM�Z�ta|t�F4��وd���)�<�7g���hju��!	�@���6�l�Q��@��/�n�Hy�);3N����
֐e�SD���X��@gc�w�sm���1�!��XR��/�3r}4�zc^r���=c��`�>��j�F�/Qʩ���B�(Y���~8a�Ӧ��ij��j���b �_.�#�O���מK�n����;�Ē�b�6�(��V��<�D"�o FJ5F��B��A f`��d^_�R��6Q�x���C�NuM�q�=:8��cn���0/��+��E^�>�/�g�%����o�T$�ۊ�)r4�r)&Ĝ�@5�%�E!=Xv��~�g�q�L9P�3X=��.�+�l��ROS�g�_�����h��E���d}���b�����Tg��9�vm
�8��Pn�T�qxj�Y¿X|��cY�H��jj9a�Q>��~��cޫA����l�Eq�ૻ)~��=ߩ�a����B\lY��M2���F�^��0�9�Q�VliN ��>��۱}c����u���D�J��e�iXqgPm[$�^�E4D�rB������8�u��H� �K0ac�t�$)�ȝ�*����v� EE���U��l9�|�g�$�k4E��9<A7�a Î��|��vc]���K��S�,Ԇ3M��=w�7ϏH��\����?�Z�2���6⩣-8-�|"�۠{��]�#1��dK��������^@H�����k�wy�KN�/�Q�xڋ>P�B�i�	��ÿD:����2तm+?�V[uz��7�O���� ��GV���+Ү|�/DjC�a&�1V���l��Z�__'�~V�s3r;4��;�j���xj�6 	�������~])E�IUӝ"�6W2�m�V[$(c��BNa�*�m���{$W�ތ.N�ɼr���U�DI̡�8�]B�c�1�T���X4�>�VŎ	��BT�~4,8�Y"a.���H/�D�ȟg�G�k:���J����_�?���E�K�,ye��8T��R��<0�#�k�h��5Ț�z��2����D�Ev�����*���r�(ϡ���k�M68:ğ�׎ ��j$�'�2<�k�(�
���l�Q]:i3�+��Ջ�a�s�~g�Agh>�Z`���I�I�!��oF�j�֕&\���p�z\��齒�~��8 ;z؅�U~�")`��c�Z����΋���/���e�Nk���@��6"$�n�=��9Q����2��3��'��Z�AĊ��b�\y�+�G�I�Ɣ�CpI<hC4G}�(�m"&$Dƺ<Q��*'�i��w�U���ͧ����m�)R0�!�<C�X���Y�wI�
�|�[�6Mx�@6AG����0ݫ�7 [x�*�/@d3� G�JH�lY5�׌?�K*�CӐ�9��\B�3h��.�,�����:6#��Y�[�9��'a������@����H=�t�+L��`�*��*r=B�Ԗ�M(QN�ͼ^$:��ЉKB:W|���zL����^f���-��4�K)v�,-4S4F�߬���]Ź E4��jPZ�R>�*5(�R4��`\�j��ViG��\�Td�g�BM��\+�/͟~������yuz��˧ C�X"-4��� o�������"�f�Y�����c��LY��ӊ����Ј*~B��E,L�ز�W��'w������V9��	38��Hس]��B�)A̝N%,=vB7��4H��Q�a2,��`�h�ô��l�l9�Ԑ|x�͔��nj|#_�ދ�9��B7��gA��~��-<u�oa���C��\����%7�9�g����zH��|ۀ.k���MO>��<��9�71A���5��Uwa4�e4�O�R�kӛ�T�v9*��( ����<�2����nI�KN0(B��|q_�2����W��)���|�q쇞�E�H�+Q���)	����+�;��[u��w@����}�NZ>���ܥ��Yzo�b|���Ô��r�\�X�N��>���93�n�?�P)<���ֵ%��X�ɣq:�ف/�R��cɆHG����Wk���l��uC�壒�aD��/��Iz����^pl
� CL����:�v�2Cm_���
�H*�l�a[#l����&�s��8��l�h8-g�=cO?�VHb��>�"�ur�x7�:�TQ�i�֤/��[�u4$y�-�#���"��~Aʷ_��У����+�,��H�N$�������h� ����KE�o89�l�2�!�8���]��s����uT0�F��K!���[� �,�\Zl &�3!�T�&a�t��L/�X(�*4[=\n�Jc�PڦsD��k>a)).�+1���f��1Û#�����J��"@�e����TŃc̌D�A�<��bkK�Y��x=��y�������8������:��0<Z<�T��J�{Ǝe��Vx�`�Pp��X�sD��i��[�,M���c���[PF�~�hZ��^�������Ĺ�W����C�KΘ������m�1�1�@v�4�dp?�U��E\�~H�K��B8�n2���Хt~�u7[K	|e�6ȼ&��~4
���pp�@�~��|#��`.�>�uG�C�xQjC��\(_����V�n9��7K�phS֮!�e0��2�`MՅLM"Ђ��o��y�%��A��Z�BY�=
O)u5�v6�����1���V���~�1Q��x�G  ��ߌ�H|h DR\��%��$�?���'2��g ��׭������1a�v3�66���)���X+�8�:χ.ȃPH;�&�Y��]K~(ͦP�f���;�0����/۸����7�FP����$��z�Vߡ�ԋz��v��/��%'���]?�w�!���i�h����3�����poID�v6]��ů�E�#���7�U`�@�it!�1.x��k�S<�3�*㗨��Wz���/�+&�^uݭ �a���
ˤ�l�5���B�tm�h�<�D`F����v�,B,��t���Q]��d<��������D�7��Ь�툲�z ���ֺ�<�c���2���M��]��G9=���V�X;1*L�o�j�9���.o�h���̸#��b�m��I����[���V���e_��6���E��'��)��|��&�<H�7x�(z�8Eq�b'��Pް�+ϩ*�����AW@f�,�=H<���D+6� ώ}�GMВ�WR�G"{#^R�ܡ�:ޥ^A��Y�.H*q~3��PF�Rn�#��Z�at!U&!""m��:ϧ���]s��]��1�.���h�Xt^e��{R��x���Dƭw��? z���́v�RU�G��=8�"�l�b$���t�w~��tĸ�߱���ZE�2��-��8�є$(�'����]��!iɻ�S%X�綹s�ZW-t�T�A(�e��1|RmA���'�Q��k�Z+�6!4��n����T���m ��imǯ��e���QD�>��)庸�Шɉa*ܬ��:Ϗ�-4F�a"���0^��^xM���&U��/L�M�� ��M��^U��
��k����dΙ��x�vmƴ�^8�!�H��PiD�맱�g�/l��R���+�6A����k���T��*��lZ�~b@�� e �YA����|_t=�,^�@��=X�O���D�5!�MT�IH9�{_��b7n/��4�rD���D��Zk`��*E&A�|�R��c��y�߁���";�� Em$�AU��*q4�z��S#��W��оƷ�`�0���Qs�9�w��۬�NTa[b��qY"Aء"�,��a�:X���M���Ch��#��~�C,�������{��¸}�=5;��3P�/,?�/�X(��K��Ԁ	oB��^EQ}m��.�x���(;�WR�R�/�B"l@Z5��NZ��N�_�cH�[oz�{��H$�E�y���"iR�Ђ�39ӫ��*�&%`��9�s��/�
�b�J�d��Lq��c!縔�����˹���*��g�Z��dX(@���C�[Q�c��}�� dˎGJ\ڊST�7L���m����������W�pdD���0|2�X2>��|a�iWH� ��h�8i3f���`��N[Θ��
	O�����PI�A���LOكs�W���SO���]���'u��29�R>�	��߁.u�eu��o�=T^�x.���q!��j5h�5�6�r;� L�؊�"�r�H`	!�Z��ѳ���i��k�0,�(^oO��s�T�Hk��zQ���������V�������sI��Cx�;A���X!���������,��j��<��Y~Lm?n��o���M�y͝��*�د��B�O!z��,�(&TB8�x֩T��<�n~w�5�~ ?.�J��`M�L̸�M<�n���Ɋ��-N�9K�<O��R*0�+RS������ ���X ��f+������\t�i�@���E�,��d|{E�B��Ѝ*��]�~��H�C�2�Lh���$�:�da|�R9`�=����v��6���������b���8�X2�5L�Y�ī/x퀟�3�C� yF�۵�{5�	8�TE�p�駰����,�j��ӯ�Y;�.j��@��j� A���a��d*�O�a�ׯ|��o��ߦ��hVƿo���/]�@�К18)�]�0�A��f�L���5���
��A�����Y�y�!����LC��^�[K�u:?@�Q�"���tX�&`i���׊~Ye���] B��g���6I�l}�4�%9\A�>0X2%�PK���gL�?��YS�D���6�{�h���v��D�&�6YF�c@炄�g��V����pl�T���`�˙UBrd���i	1�i��~קd�1��8
a��~(�E�f������3��{6-��ha�(�-'V�f�'�%̾����й8a�
$?v�ج��ֱ%�T=���Za����0ػ��pk�#�0��^��Pf�`�f�|_�T�x��g��J��J������ӡ_�!�0�%�v�`9W_+4� �X&c%GI<��<+���!���I_]�A�.��Tz�ފ;?���^k�x��]�3�����DQ3����B��MM'G�D��
#�<WB��Ͼ���SL~�O\3��!0)&�������er��F�ؼz�u~Ύ����~��sJ���Piz&��,����F���=t�jo/��7`H��V�vTp���C�K�K== �C�P�eG�X2����Zs �W<��N��6&���X<l3�����<4d��1� �8 �F9�y�x���	n&D=x�T2S�y�ɽl�1�[GR����g�(fe}(o��$FQ�=��co	��,x��X���G��
��P�>[V��w��RS^!�t�,>���Iҿ�U��P4M02Z��Һʋ(�=&��I y�.Ϛ��ŭṢ_�O�Lb��ʨ �vۇR󔾒������J�sp�3�ӤI����ׂ�oݜ�Y�B�Jw(j
��|����a���0>� s�z���������q�=Y�A��o@���|��I$"6f?px���h�j��M�C�;Ȁ^�+҆������c/b	�p)2�e� <p��\�J���>�r�QKU#���NHU�U7�kX�ܴ�����F�:�Ԡ/�>R���˳���_q�U�������s�h�Ř.IJ��X�#�|���!���&T���g+���*o�[���?����ޑ�4 �}H�'�)`�moV�`x"�,n���������$�l�$Ă�v�( �L(�$�s��uQ�y$V��i���ȇ+Y�<|#,I�\��΄�0=�
�P�'CI��M�D�����hr"u�����i����o��Ի0W���ޫHE�{�;K�(A<l.��G*�
=Bc/6o���LQ�ٔ�S�π�!�E��!��}�j�T�ǝ&5�AE}��u���}*+������j��.M)j���e�|�}<S/ɒQם��#p��3�?v��EK��/��O}
|�3:�y���u�W��ƨs��\�����1����À��2�W��h:΍{��]����	s`�Ջ��x�ݨ��:�/�g�5�f7����W�_Iu�7�♵�c�8�ò
��+ѥ;��<�$�TǄNX��l�@�4U&����^��QQ��n�~�k���� +���|h�x�j9:�ԺH�^x��#��ss�:�����<k"&~��p,c������Q��2�_r��K!ߍ�������vz �)_��a�a�x��NV�IyC
��芥W6�PM1���E�=K��,jLu�R��ȸVp~���O�~(��~�VBe�ˤ�|��W�#G��#��K��Y.�6���>����O��]�e�������������}�c0�;�	���S�!�w�N���{B�z%��R)�&a�I? a�/�@���gh����R+�x7�OO��.Gԙj����W�>O&�\���(��-�M>�Qs�~(vwC��1
LC�k�O�P�]E�a>f��3�Z���G�H�p�K-=�*��+��a��5���K}��������by��`����_2�,���C*�Y4a�3]��s�a�Wl|n�?�Q�����]�$�s�
[�#����C-�E���� �����O��� :c����֤#\4 ��}�S���y������\��(L�H���&$ƙ�vg����n0���(3dr���?U~�Ez7f;R{&�'OY��k*}��s%����OE��K��N��(X�:�%�%��`���r�)_f����?���:j����������]��[�=��:ES+{��}�-zֱ)�ι���$�eg",�$>���4��U�K�5��L���_8G�4	���)J1��m;���%z�a�y��r� �i{b�d }h�C�����ѭ}M�ڠ4 �(^P��b�a�L�lg҂��>��׿�FZx�1#`j��s-8L�4ŤY�ꦐW�d,�cެ�7w���K��b�T͆V��&�{JFr��&�_�����IqǇƲF���ᣂY�{[��5"h9���)���.�éaq���	g������b��D�2`<��Tě�2�^�w~��,,��&�˒�����r�V��Ro�L�)�k�����F	��`��ۺ��uN"�x������4���~`��(�F^�L�fǒ+)#����<�8�~�.0�.Z3@�/)+��SU�n��=g���E.+!����ԬL�z|3l��\A>pr��M?���i�KN7E�=;fH"؄;5B��GM�^4>JzX0ԫ��q�~�JLO��A�0�_(.��*C�@��,���@�>j��D��X�G݊h�L��#��~���󮲔�Y�� �F�~ျ����q3�D�lꡊ�
�(�X��ܙFEO�cOmEV sҿ,���k%66�g !�7�������'9!a7?S�H�YӼ�P��n!� �Uv{^�P-�n�Sp9���Q���Tx���W�
�.3���d�u&�E�`n%�?%sp0T��=|s��쏂������h��^�=e���C�z����q��� c%���=���_����mڌ�J/�#�/&[aߘ��N�	y��Sy>��+�-fJF�`$w�7Z� ���4����������b��o�d!x�΂�	��U���5���>g���6� @�)�:�N(Z�r����b\�*���+[<��B��*�6�����y���~�W>d�E� i����h]L�X�Ϻ|��
���D�G_�$�8�x=�m�Տ��c|h�z�v���ˁo�����A�Aa
�܋ڍ�	\��U�
�#��J��ǔ�Wd����k�����!�xYQڃ��vC���ye  �Ǖr�VK�Jx.&��x-��PD;g�s�_����T��!?�i��{��N)�{���tͻ����Q�Ȗ��t#���O�~�퟽�6�W��ڵk���n]���szr�猂}`�d�	$k��b�DT�"����fo<��A#��I��x�:� D39?(�3L����T2���q��<ɣ|������r�!o���z��J��>$�0���+o8 �����Sk9��׉���H(F� xRb�h� |��&J��dF��5z]�2�![	��`�L�q���`����F�P(��'%)��('m�Ĳ^�]�NO%��Wf�  @ IDATZ��^�����vw�7VĻ_-᭠�Oo4��Є�oXSX����/ ��fX�67��z��,	
RM����`(`��eƶSs�v�ǈ����ݩ�PPԛ����-���|��tA*�?zpOt���������~�e7�ãC`w��&�۬E�ljX8������|:�>#������}ϒƆ��������TI�=�۞P��D��g�W�ҝ*3��^�����7���{�w
�
��{�K~�([J�}��c5NV6�z6��,}_$�Oর,r��Mx]D�H	�@�8��?)_u�=��xk{�N8��o�o�ل{�B�28 z-8Q���/Oq۲���$ˊ�d&%$��QC�U�	1�$@��4�T�d$�Sʤڨ�z#�$�I&�g�ُ�Cc�b��l&|#�y|	���~o(�����$���0j:B ��T��t�E,bH�x�����ˏ~�#���װ�	�������"H�=͊G�2x�ǌ��l_<��L��/X�����v�X5���c��وT�ZE���rQ|�2D�|��G�N�=��@l`���E�2+�]�-DQ��g>�eK���5T]@RFcRY5�B,H�)��`��	(q5�u�G�5,#T���P&q�ś������z�Mj��|A��|2��)Ɠ��"��~���	�	�v��f.߁�jNlܝj�_Ѱq�09��x���%��	�s,G�V���jPO�IY�$3G�l�����	�èY�j�����3�g���-��~�M�d�� ����|P8�w�?�E�G�3���ǻ�>=.�BO&����Pv��{�@��	?"��xb���9Ax�SH��V 9J��s3��di��%�����f��NO��tZ$�z�v��I���N_�p��G�˦���{�@�+��خ���o.�/-�����[?�	yS]���*<�� ��q�c�MKP�,.`�#�, �K�!.�'������Q��7Fv��I$M2�$w#�L���ǋS��:��8�6������Z�6�ڇ��U�R�D����*��6�� �
������D"����o�܈ F���������Z�<�����j�}��O��A`SE h8ɷZ�O����őLfڵ:��h2bn@Wp� ��.���tt	��Ӈ��2����r�v��3�H�Ue�O$D	r��-�����~�ӦtwF�@o�(ܝH؉(Ep�h�%��JM���7n�-��4�`n�����nj~�vr!�2Ġb�utnd�Q&��ƃ�
P���Ns<�0MZu���i���Z�lsx�7����X�
��<��qI�'\�O�r��B�c�OI�9�+� +��O�7��0r�$9�r��-!k]=��H�Il��=�7;�h��G:�C%��^^ݾ������ɒ���Yβ�񈸾6��]�얫�n(���~�{0�!�L��|�7��3��,v���'j< ��������o���?8�!�����RҤ��.�; *x[XQ�re���CBj���	l@tQb�ג�O�Gf	1�];� Ҩ7���ccQޅ���v$q"ŋIp��o`a��r��Gz�e�����a�4,<�-h��� Eݱ��Վ
��9��#��X�ވ8�} 儒�RI����������OJ%����})cۯd�3���%e� y3ӫX>�*Ճ����w�|���!n2���1*��8:öfzD����v,�h"JnM"�"�gH-�O��D�W��T.��YU�D����6}�$���a0j��qʝ��H,ݤ�"aA��Zcp�W�Y��I�I怆p7�`�[�p<���v�Qŷ�{o=��`�5��<�3@i>�FT��W	�xak�8I���h�r��_�J$4�X&\h9K�A,�{ZÚS�8t�\�OCj;�!�*��Z&{\8'��X�<ll#ˢ��j����IPW��Ï�#�7��9=:bmL�&�N�"�
���Y2���ڡ3�ŕ�Ò��E2D��rL&'Ǹ?�7���a��5LM\���{)lA��!Z2X�#��]8	f5BL���jakg� C�8�U�p�W�	��8�v���<����4x�M������4�W�%1������8g�?�����`��m��b�(��%�l���e��|߼y��W_%�����������v���I��05u�S>�����/���ē��E��-V+]�T��j�'�,�8h�)��� �
� �A�&�M��n[d�xL��z���,A�H��>�o�`FY_4��'��ښ嘭gsx\��EoAP�`�A<��r�*14GL968^��p����voow�r��X���E\���)5� F��$�'��r,��Q$�麬�o8|(�"��Pј��y�����yo`ﻚ�!{��90�M�p"H1��tA�O��$&��ge�GC w�j�t� �:�N�P���j�d��&����L�g���fҜ ����dב� �X��Z��[k�'�#���l��P�pR`MЍB�:��k��Pp�mS�\�,F��㲰�1����|� �KY=�U�������Q��3M��*�(��e���NNN�ݿ� �J���%<_�d{����B3g�ɘ����1�!��s}h6Z��?���<@��)n
�Kܤ�a'��F �����[	K��p�J�8(��'���I,t���c�?<:�������e���$z�8�O2���#��F�TB�D����i�L��/������L?ML��z��i������v�.�����j�w&�{R�b�`��R!uek���=�O��o:8GNcS&�}>�=1.�߀;�+0"��c�<��d��Ą������t��(8����s�y�U�����a�B�
N�0*�&I�78E�z��dG2� ��vr-�����7��*��*�h0D�"�@�Ihv{s���\�YDx�!����PǥϮE-ʐ��6�ϊ��b�s�Ǉ��N�~��<�B6Ʃ�(�:��X���bI�Nz�N�D"�	�Ҭ�|��o��ή���Z"w�ߢ���Q�sk\,b�����5ㇹ!ڣ��YP��&5\2�]y��#1�PBp8�`�F�\ ��
V�$Ж��X�'Vk��Btp#LCI�D$�9��Fa$I2�泵x*Dɕt�5��O�	���ǅ��zj�IS�B�EEM�c�ܯ�n`�ω�r�(��z�utJ�<�!%=�n�eٔa��Z__G��Wq��M�3�IL�g�s��l2�uM�V&`���⊞���L5���/߼^��O1�0��`�q!��81�R���C��rY�A�,H̝�"$�7���Rm�ӗ���n��L&~��!���H���< P3�0��P��n����~x�����剆/m�L=zgB��k�:�>zH� >��Y)bV�;$��iQ�8�Q�-�Gtqͫ}�ʪX�H��V.J� 2��x��kW���l�啟�����u�����Ee��~0����b�׾���^����%0e�ݥ��=��D���0'}Gԍ΋v��JE*P�ܔ� [CZ�?�����;"�6��+�Z��W�]#��'?{a ���t�RQ@Ȉ4��d�����ē�.�2jI�lM�Xi�z�,I� C�v o� �K�x�7���q�C��u�j��j|�X[�*�+ky*{olo0X�G�db������������'�h�T���ީ�8����B�/6j�#��8��=�}!>o�ǝp�Yĩ������ vn\���zppH�D�Z��d��"q�'�����/�&�8����?����^�} �E�%dؤ��#�j�����&�t,����5�h����|?9N�2YD��*���±=�)�Z-g�
4�v���O]Z�8�(���f� \��@j�����{�~���]{��7i�3�3�X��+��ڠn�����oo����c�@�B��6I,�S��'�ތ8���ߺ��D�:���_�b4���[x��ve�e7�Uь4�xlĿ"�"k�=<R����i8�� �X0�9BFr��Z�!%�k��
2�|�X��d�])M6z�j4�A.��m��L�|�~���r�^� ��}�����8C�=ϵ5���(���gC`=(��I�hZA>����Q��)���W�7+�F�e��]�vj�w�m�c'��Q��=w�5z��,�V;��o�R
�E��\&U<W�_���t���<�]sO�k������=�� f&�z���pP�t��y���p�;w�?m7�8�!ƌ�ǒ ��I~����d����GH()����YQ��TPƊA?V#����^Щڸ�}��S=\�R�-�2�dRY� �H$ ��3�"m _8K�&��$4I�U�#�?����k���a�Ͻ>��Ӹ��qe��߿b���#�Y1d(�Je~�t��I�%���Տ������J��fD��a���̟�r�45�\��JJ���ш�� ߼|	���띎�#�@KD#��4��St G �n{s�!��E<g��Qq���p�
~'s�S���\-�/�r��-��xf^���^q�rј9�]���j���]tL�.��r>:9z��^����G�$z�W(�b^�����Y�|Ʃ�B-X����E��5<��xX�h��$S˥�K'\iS�|�x�����ε�ˡdAL�N+e|@��[Wo3ݬ��~LF>�6	������@�)A~���^~;o��G*�%ӕbi��T����ta��E0'�j(#�I�n��$T��-�C�=����X@eg\� Bt\��-�m]]e��/x�t	�ף��!D�t����B^�@����|&s���n�p����?���%l=x���n
�6�Tb`����s�<�ee>/>��7 ��$��g�0e05�:@)���G͉;`9*�p��fgBo�x��\��%�DH(-<G�@l���[Wp
4�?�i�t���I�G��=5��c���a��GPk��F$Fg<��<[3�J�� ѓ\�niv���7�n�V�}�����l��+�?&?�~�+�s_U�*���k�����K̋�d�"G���� )�J�j=�E�FH�+��N�C(���yi}�}x
�����/M,�z�1Bʝ&�0�;�-��R���;����( ����/ܾ�����.�|��Cn_��<9:�r�����@i~ݑ��M\k�]#��`x@���Z��
�8���>��l�x8a\l�̤0�W�����!ȇ�#�mټ�i�=���&<P�Qls�٥O����
��ñ��������/�JDd!mX��A�TR���)0B�1G������J��0��[����Mng�&�lK�X2��A�.��Q�at*��Gcf����
j7!�]�N�*x-�Ô����y񅛷._#e=+P�&]: C*-X��<�n2���6�{��F6�����I" v (=)��7ƃ*W��i��6�E���c�_5�ˎ�����c�eO����W�Ll����i	����>�2�8�:I��j��� 炴�ΠOB!�]B�"������QW�U�U�F�3��|	�-Nd����������Q���N���ǃ|N���v��= �T��/A[��t������ƭ���x���������&|ɮ��Exܭf��2ґ�{<�q�vA����P .R�?�W� ����2r��j�PE.�����꛱XQh�t���s�V��ӟ������
$��F��ċ���u/���Tp�+�C�5%x��d�SD��{ {����GgЀfػ��7N<%��C���%�6
�&�f�f�g?��I\"��2w<��f���s� ���nఠ$N\�~yJ�P8�,D�b3�t���}s��f&�o�͑z��^�#�9�0J
�f��&�bpZ%;�q�'J�ma��ε�7)7Ԣ�=��aPvF�%F�fY�a������1��)� �=�1��/���C$�)��/ˌ'�Ht�˱�p�/K��Uܭ'�Y��8�V���7ZX<d��X�6������/鱓)9y�j�4��E� @�ǋ��vi�!�h��$��CBx~�'s����$܎H7�8<��ē.ju p=ڃ�,o���r7Kj�"�W��E⁫qGj�&��p�(���� X�����0�]��n<���~��Kr�,��B��ǯ�c���i�W���O�N��9.1Ϡo�p32� �<���� ~9H�)�@H_T%��c�	uJ��X�<�������R^�E�S��7j�{�'�&Ҁ� ��MFG���#�i�ʽp��v�+�q�"�+Wn\�
'��!ψ�E1�d.��R��D�!��#�՜M���-��7#����ݾ�ie�(�s��E�JŘ{�0'P�*T��s�+O���O�Ù2N���4��H,�@i!2�l�N��ȑ0ևx"`ܵ��z���]
����JED�̺z��gd!YVr-kyu
��T����x������
S��B����>H��F��iy����ŷg>c�vQ1���3Xu�p+�">�M��Z�o5O�޾1-ػ�H!��[�ګ�h���+�p:��/�:��;y�!7J�3���2Y;|�;�1W<�{������ݨ� �]�_�C�uNj��G���R�^��χ����� ����fG&���ɨ�e�Xz�5J4�=٭xk��
��pG�N�$F�bU��M�g����d��/��_@6V�E��z["�ȑ�K������,>�|"�X�<���p$��=��a9��*&�����d0E����ްt\ �G�z��㒌F�ɕ7^�
�<�-[�<����n|,���Y��E7`�(��K��1k"�e"q���f�,�d�x����K����#�~�����z�N<c����&�	��܏�xv0���/ŏM
�`���=�Pi6'�o��o|�G�Qf��mIq^"�UHk	iB\S��$܀j��r��rLeJ�ۺ/��!,�5�����K���x3j�!���}����|jC\�{�����%�M�j�,+�1�$���a�nQ�|R�<oMƼgg�h�$){ĸז�z���k�Q��j2F�*;(�8�0����;���ɦ��e��ᄭ� �}tnIvR,7�|�S�l;.yt� Q�4���YE�@)J�sF8H��
�4ˣ���u��N����2��pY�2�}�o����/]B��2EwW�A����!����ߜ?�u��t�����Q;)R3�tnvstWb���&����:�hY������&O����ޞ�J�ð��h4�� h ��\�B��v�Z�!�t����a��������?9��w-?9���Ö̰LR$E��������2�_��Ϳ��N�����v)���P�NUVVVVVVVV�	��K�d�اϜ6Xo>}Ɓ��6�*��8�R�����׿��_��y�[q{)!�|�7���{����L��ߩ(����f8���o���-�DS�\�WX�_��6+����8��1b�M#�4>6���[Ώ�cǤN��C���Hgp/���u-�;D��{R}��J�5��a)#�-�^����-����p�d�Du�(�{��O1>u2)-$nP��3��dk���o����7V��M�֐U�&'�Y��q�j���[�!þ��?����Ye�	T�ሿ|t���w��z���y�����|�����~x�6qn[kT<��������+<���Tn�x��B/t���t|�XǶ/3��G�����_��3ܟj���}�\O�?�#�om�{�|��>��_����l���1N2� �}�3[����O���������~���<�����������_|���U�\�·��?���_�lbww���c��R���v�9�vb���/���68s��t���Y��)�b��-g���r�������ERF��N�1��n���0��Y�x25����K���j�0�-��3m�=YH`�k-�����t�SR鋕ɲܥ�����uL�P��(�4Ͳ��i�AV$�\�zI`����7�\d�PEv�-�L��,).�_�����#(?���_~����������b���S8`yk+�������^f4�ٟ�F_=��k��W.]�u綊8�1|�tΜu��i^�lޖ���`3UЍLC�ƣL��Iy3rqf:������w4%n�a5"��[s�Tx�|��_�3���'W._t����Yc��./иj��W� ѯ߼�ǚ_��>��������������7���K\=}��M���������CN}�)/w_�;>X�M.��˧Oy�ٴ���nA�ND.(��>*�zV��y��o�e������ӟi|��g_Xd.w��������������f�-�T%D���������Ũ��b~�#�՚�����T��z*�b�=�<E�����ʗ���{z��]��OflŠ0t���o�8�s#�g_I^�lm|��O]7������/~�����ROٸ�p��);�>�y��?�l�X:y��3Ow=p��K��Xl+·�?�|�e�B��阴�Q{oI�٭���K��q�������
��xx��c�(�����֨������g��0Swu����S�Ǒeg��f�|dz�횦��_<���G�q�����K����{��iL�X �<������1�G�e9s�����L<P����`�&>oܸ�6���z�陳g�<��|�B�w��u�C��L�*X��w�?-�T>�|}��M��8Ǌ�4���?��-��1��@�c�N�i�:|�&�<�|$n�p���	.֫����T�N�����i+O���[s�,��|���|��"�"c���!����w���+d����⋓G�9���G���z|�cR/^����׾�����;$����B���.mx�[��ձihYj���m3����l<�m6�͡�wD:�׈��q�	��$<v^����On�vфc�j:����w�HhVK=������p������[w8������7?��缜=~�9e���:���G�^���f��������M������J�s�D�ܵo��.�U\�������u	G��f��'��(E2�Z��b�f�	�@��E�u&�� _4Z}�l¿]��Oz<\Y�b�CM�p������ 1�	Ii^-λ��1t�]�X������N�ԐZ�8�o>�{a(�A��f����S�d��O�o��@�E��m��Q��~��gOl��y��<;�W��s��Ű�p`i����{��ᬷŕ%�@7 � *g��ﭝ�x�֍�l�X��zq�;W�>��� �Z���֏�ӜJO<[�xL�X�o�
���R��q�Y�����:pT�]�q�d�1D�Aگ?D���(�� �?J��!�����g/����~�ז��u�.+!맕9j�+J�yhM[O6�srf ��;6��y���kq�.�x�r[˂�w�я����ާߵm����G�����~ĳ��)j��ׯ�����g�d�V�jЇ��ڪ��ۮɎs
�ͳN�����Dsև��FZ�vbs6�@�q�Z(�ѵs�R�co���\�}��kʹI�ʇj&oCY��a*����q�?�n�y�_�\�lO�3HH��C��� Ϳ��E�ybϏi%Y�������|��_w���s�����CNaS��n@	�;����/κ� uG�|����7��xJ���o�ʤ���v(��>����O\��C�ZB�1G'�v��i,U�3n�ުs���;�1��O:��%�U�����Ӑ�r�=H.�������;���O7�ɰ���G�w��o�G��pr����;xvq�ң�QVO��S�6v�f�J����\a��st?��\n��&6T���~����fA��Dh|s�M�,d�C�������PO��Z�5)�v�
�W�|m_�>�i���1|Nz��f���]ʲ�İ3�`�eH�P�fPů�u��]27�9>?�|x繓 �b��;�f��Hc��0'P~b���1�l�68�ay��nz;��w�ĸ������آ���d;G�6�GKK[���幏����6�;�u{Ӂ�ny�dz�ظoQ��9i;����u|}����Y����eLp�`�q�7=u������/o:����>���(4�F���n\\s�0tg͓�l�W�^C>	�TF&}�,F臏�3T�����>0"���#V�^U�9�W	�J��@�h�CAN�Y:�����%�%sy������#��hu���;���w��[*�^]9�u�nc��3*�xȚ�W
Y�'K˔�kW�"{����Ǐu�������!���e��� �H��>g@B�xR?��p6�K-w��w�C��_��Y�>���$ J}���@�u[4j��Y��CF 6�8!��D4��Ⅎ6K���Ob	|	^�l<�����}�M��{�����H-Wb��P�P�ѭ�ܿ���k�Iǧ��������8��Ń;��b!�d4���yV8*����Ο������?���G\d�-�D�m*�X�3?bHd�snF�+4+�ӯ"Hzu�p�����l�ν���IvY��o)�/� `�8q�p9'�oRiƯ��mí��Q3�+��W]���u�Lݜ�},T��������L�ݐ���l.6r����mu����R��:*�0��o��C���8�rup�ۑ���;Ξ]�x���i��ԝ,F�}7O9/tk?�ɄV�dbF�x/�bB�nk� ����a�R"L��	��q��r�����OCQ�I�`�����Y�1��R����=@��/+ǲȳ��cG���G.���Y�KF���JE樆��&sEx�5s�7�R ���B�l��?��ثy��7�V�ѐs�(�/vm4#У1�K��帺����]��-m?z��G��G�<��υ�n2�[p��h�0w[�VѨ�	<y�1����GcbeYDuDx�--�0h��!��R����br�X���l0��8�	<Bm	Z⃡c�H,s:u�<3[�ӟ�����!�#���y'%P�c�O0o��ogu�x�4�>�L�]�pQS*áD8[K(PJ[h�Cń�\>��x�*��?����S��6*F���2}�2��� �*����>V>�J�W+��i4bŧ�5<�5���ע�ņl>dp5���[8 p�ذB�h�Y�2W�[����M~ DZ�SD7e���L�(G�Ӗ�L��ٜ���b̨����`��c��o�r_�r�,7#�{�>8����?��o��؋�Э�~ɒ/\8ϵ �O;��w>��Ɠ'])�r�D�d��Í'3� a|Q�º�����8|�5�I�/H<�Y��?ۈ�cC_<)�������L����J�ԙ]]�WW��2��悀���g"Ƴ��V_�����cwr!ehq�����W���jn�0k�	�rh6��z�J.��Ǒy��� 6;����n[/w9fݿw��'�����_c`8�H7�sFM�?_9e��j171�>&K�����7�?<ǃ��%���^�,G��e�-��$�Ď�7�s�"x:�z�9��!'VjQ���
&�G�<4I4vE$Ic݇�g\�[��7�'VI�>��r�}�!����z�fu�p�Kgiq�A�O���K��XILf�!n�[�)�2����L���V�v�x]^t��Z���M�J^�T#":�wV�)j�Vk*����,�}ŌK�4�s�]s$��R���5I���4�1�-�4o��|��z�B�~]��s^�V�,!�r����1�Z�����s��<���{~�4R�je`��<N�Z1^A��_��3MPpә��q\��]s7n/-ԋ�H-�Q"A��������,�&KM�%2#4j�_���Ġ��g�M�=���؎�˒`z���0��8:��ٵ���g�n_>c�c6>���ŗG��>x��g?�e>Ї01s��Ѹ&>;�{����X��U�"*�D�7�������&�Wʕ=�V�yf�}^���'*0�N��d�����W9:cpd`H��r�� u�|�_39<)��_,<QD�+��i��m�!Y�o��X�+����1�3E|�;�c�1�_<��G�e�JL���=��v�`����u��`<�+*�d�Ї��|����y�8�w͠�r�?B}!ݘ�� ���r m�_��;�r,y�!������-�]����f9��E���lS�vr®�O�W��!�c�(��4ǘ��	�R�\���/�(=�q���ͧ^n�}�������{�hg���۝�M��=�h+<�ay�no>��;�!��1PB�\~�L�葍
%�D&6���ݻz =#D����BR�;��`2�{r���Na1R��_���e�93��R��E��~h��q [���P �C���p�X�@��k$��\��NVp
ø�����_�H�G����;�7_^�gO��Z'�>l��!��&ξ�urq�B�-ߴ#^V�c�7��[� �<���S�_I0HfD
���Gd郲�T�eU�3����T��`��6f,�c��������yD����r$@�/��>A�����g����Ҡ�_#uNw�ܹ��'�����i�4B`�͌�4GJ��r�����/��~J[�K+N�h��oܰz�t%;q�n���Ņ����h�-N��5�O��X*Fv��I�F0��#n�-ò��fBb+��i�8e"V����C��gP��?a�g�*��R�s��?c&�˾t����ɖjaD�c��SC��X�Ƽ�X�՗_���q�&j���n(���3;��{t��~�A��̞y�Q0����i�L����e�����e���o*H��Dw��Y��t�q�#����~c6�yp��P1;�FaҠ�eSƌ2���~yS<���s�����i8��D�7wo?�z.���f�ߪ0Mp̤��ө>z�cD;kik��$-���Zo���Sg���ոWk�E�^�<�\����3�Umzr@��n-���8_^z@�C:�5�O�FaV�S��ƥ+�����VGz>]�+�����8� �Ȕ�;.�Ȏ5)}Cy�<{��Pn�Kd&wd����8��x�:��֭K6� E,������V��|�.�)���Gq|�ݻ4i����sz�>�h]��q�#��bүv`��fĎx�!_��9U(U�k9��di_�x�� ?�c���~,�E2ȓ��
�Fx]�FQ�G����c�#
������x祶��/��ƍ��j`U�����a���!M�� ���QD�����"��!�m�q���e�r A����l�@�j���?eD���fw�F	��|������>P#bLTI�R'��q^�����C����Ej�.T�#� �'`��R^%��Uu5x3������Qk�ֶ�h� z2-Qo�v�2�������4dX$�j><�F�0';C�p_��8
���,ǖ��_=qu�Sw�Ա�;q���;O���8{��)���|�"�dy:�ǿ^'>u}Z��|���6ȹ� o�k$��ɺ3��R3HO*�Ր��.���׎O%\�cq܈e���p��Ot	5
�*��c�|���[v��:�@���6��w��e���C��fXذ��S�C��5O���gw�9���b ��p�_x�7�a�Nki@��n&ź,�(��E+���d���(�w1q��~��8��X;4�b'ۚܾ}[��z)���׮�
�ʰ������_��:u���1��cD>.����>{���
�
|�y��3�"��Ϭ�w�Ύ��u��|���+��c5���X��#����9���v��s�S�޻u�/�kC���,���I��	9�?{�\ܽ���I�������C̲�[>�q�e"�MO����s�ݞ�.�� ������kn5mܬ}M+-�h�#K��$��͓��B� &�*��V�0"�ʍ���ʀ'j��.h���<�e��yl�ۼdU����D��@%'u��h[���?M��R�B���61��N�+�(
r�"lh�Wl
m�ސU/t:��5x鵱�Tv@!G��>}���	٘�`'��C��C�j\��fS����������fNbx)�'��f�Ip6y��ERӕ%�I���f"���9k��H�F}|*��sg�'�0x��♳�<�UA�H=� slͱ��r�dh·]8�����ʚ)�>���쿠c�� �\賻�[~����G�Mw\L���|���
N��ǟ8๛���,.�Bκ�H�Vv����p����g[q`#����� �9[�W�P��p��M���!i��s%��b�����.q���0x
�/B���1h߽��� ������-L���5�C��0���/Q��Hm�s�/y�/*.JGq�π4��Kod�޸A�q�9����]�d8^8d6�1@GO#�'}�	�aī+J>��ܔ?��#�>�iƩ��/\��^O��1�s�ώ�8���;~�޿��:��u6�p��n� d��u=Dv��N�w�	��V��7���d�	��ܡtH���I�hE����dh��s�jl�� B���|���������������c�rb��g�jJ�|�lx�It����T��&��?��N�D�����?���k�n}~�ʕ���;U�T՘	����_jK�7��,l�>p���k�H?�"�<�n�4�B��͚�v�P8�y���jg�?��)��eMc�k�501vQ���x����M+�_?���ajj���{v��fCpҊ��+f0��������$L���Y��*��y���{��O2��`�i��y�;����Ӯ#]'���]�D��1j�5�[1O#G����ur��M���@+ݸ���P�����e��K��u����C�w��ܦsK��w��->�^8�sz�����N-��?��?8����o�����Ofp������������۸P�6��&�'q$s9S�Ϯ}����3���{wnx���?��������;�����7�7wcB(!ί�P�Im.fڰBl�/�x���֗���������_|}�������ș���nڰ���M��A���;��y�W�m���6^��'���6��XZ�j��@�~�X=����������'⛎Ybu�+G�)��9�8h��#�5����-��\p������틢)��R�Ȥ�m��z��'W֮]���-������D�$L�w�?�~Ƹi���܁:�t��Ɔ$s����d��;aMB���l�O1*ѭ|eN�~�2m����YX�&W�=��l�1����������7>�Χ,��o~�կ�{?��'�~��g��a�`�-ݪh6�[���-��QIۇ�|��D/��X������,ݯ����-T���WqSe2U����+�'�?.��Q�����2�nZU�|M�0��;--Cjn�GHj,�81�X�'ˤh0q!��r_���
u'�M��F|jp�#�<�k�?-{�lhE  @߿��$�����W��?]]u�'���G�?�X��Wa�s1�6y�q�x�p�@H;O�P9&��'����_)��~� ��t�杽�~n�Cϓo�^8�n*s��_9!������ܿv���/�v����{�9���S�1��>���)SN.pi(
�3���y|�+�׷����_�����/ܾq��K[U-C�i(B�몔�3G������}|�˯���c������;p�?�3�������V !Wʏ�'t�B��=�/�w���;g?���5��o�s_�qg 3�{P�vO���]�T�4��wg�Z
jN1�1C,}Ţ<�grH��ߐ-�Po�#���*����C�t�3��j'�
���{{8�).�A�#\���^���E��?�k&� �*q�~,��
A PF�=�|�	�1����̋)�ZZ�9Ehc�,�5�:~|��͛n������%rg�����x�����ͥ;n!�x�̥�?��z���ܫ|��3ۛ  @ IDAT�7�\����[_y��O?���K�{���7�����_߾m�).�&|��FL��0��V��O>������x������)���R3�/]�q����ݸq{��D�ϭ��
�'XƳ��qh��gv�i�׎`t8n[:||g��Y��8;9,$!I��ݤֺ������ڰ=�!����B��wl�"�\bk����0������f�	�Ce��V�Fҳ�}��;wn_�t�]�~�;�Tj�� ���Uո���o�����%f�
���8�Vvޟ���7��ʝ�Q]�����|��҈j
T7)�Y&B�*O�,'�9��#��m<��������_X��6$S�S�L��E3��t������8�ѓg�6ӛ�ȏ�9#P{>ֽؿ��8*�Ρ�R=��Z|��������o�v]{�D���uc��>�������C�z�U]�������O���c�VM~�)�1�=��q��ϡF�\]U5~$�ى�F)�1]˱���W#����/6�33G�mU��Q-����8|ы��D�*z�_�Z 	���P�oL����U����h�c9)�hn��`!��H�iL�5}(2�\'&�^T����4`5:w�M4T!�g��@v�Zx��Δ��V�Í�?�|�|�1<��Z���$���cq�K�{"CA��"jX����[]�'���O��#:>ͣWTX�ݗ_~� F��f�4E��f9N 06�y�TK�3�9�>i���a��o�����@m�w��6�E@\X:*�Ml��X<b�s�I�o,�4[b5��l�����!J�9I�[��1�S,mD�tf���UK{N4����{}Zl� Am��4|Զ⠪����W)��M߿x���C�Z/�9ꤛ
Xy�<�{��;�:��굫�>qZ3@R:�����`�����(���X[s4���)�z����u���|է���w�����������	�C�/*rRZ�� ��(<�cY�o<Jj�I�⯤�h����ZE�de�!-ࡩ��~��zȐ����B+G�Q$%������Z�x)'��4��pl��S��>s�5�ͱP�CY=�q�h�u̓{$�����H1�1��AF��u�>f� ��� �)S�?�X�F9q�zmYΦs�9��eQy�g�a�0����m�C�#	-I����C����k��*����[��;�X�F|�����}��:|(�U4�c��ҕ+�C�ȝ��[�ˈ)��٘��/
M��v�Ѡ��-�DW���	ˌ��>C��Pԏ�܋*}��^剢�݆�fO�{yb	�*��V��X���݀W��n�+S�T�5��o�� ��T>6�jo����\��8I�
��dw��=�~�(0a�H���g����}4��p����������@a���X�6~cXS�[�g�NR�v6��dv��a��N�d��q�sᐘ���z�"=�BK��
=v�d������H���Y
�V�Yu5���Ɯ`�.�8b����\1��$ߋ[?}�ܺ�^��B�2`۫�庣`��7_��/)3Nt���d�!w/�^����l��0M:F�@ͯ�$�"�҈�3>���S~��>°>��^�"P;���ȒE��GwD���CkL.rICa(��3c�|�S����<G�__'T�l;7�;q����U%�A�I�A�B��xx�\��n��-D[M���k7�4��B�V�"��6V��u-s8G=s`�5 �"h���q�ܣ�R��OXz�0���9�)�R$jR���J���L~c>�<δ��u��Xg��{'��%V&S=F�hW%�p9 �G��rz)�daЕKc�^a��G����L��1(I��ҍS���T3*�L�ͣ��h��f��^�Zv�bO��pƓ8	�|V/�K���W�ȇL�N~'�1����x���{��A�������HC��1�Yp�!���2�8s�i�e�4R�nm]s#J0�a@�нE�Y
�
���o��F��aXpj������D�����k�U�E0����+�|���a�	_�9e $))Gq%y}bZ�2.,-�w��}�}�WIݖ���B�'"=�q0y�˽$Up�y��%��RS�$Q�7��` N-2�������_De�&(�����A|�
�1���'���t���u#��-��.���!���o��;��Xg�O��]�
�U�F-�o=hQ�'\&n6����.���q^�bWm�gֱ��ggN�Uj�!?� W�19��E�b^+p��������(1�{��	4I�i5 YK�P �8ah���р�&�E��iY=���t��߉���U�M<n�R�1gk�h�:-��@c��CBi����)��p���
�81F��Lħ��.!����f�i��T>����ܭ	'�2��������W7�Cг�|���iv��@R�4BA8��(a|O������oK�W�Z#1O�Qn�!�ŧ&	�y�O��	�ن*h�R���TPX��������E��e���(�Q���?S����0��s\L��UKQ2ԉ�X� ��m��u���lET7:u0�[��:v���lq�~]�o��\�Ŝ�m˝n˒&�`��H�v�P)c�c�I�d�,Nܻu��&��?��C���N}���Z0��[�+
�!�1�EVkK��cY��8!A�2�+`�����CUů X_ۮ��W=9�H�3T�5�A�d�yqQ�+&E�6Ji�Q�Jm2_+��k	�+��3��3�?M���ڶiA%�e̴�PU�4��.2�W�*��tHg����׏K��vf���U%��,{R)Q���c"�ʀ[ �(����iNMCyU��5�Z�P@����7	�8:Qr'��5۱a�{Ԣ����EA�s4���kO�
W��L��1đŃu�
�L��|�a2b���I=���RLPPS�:$�݈�P�Ż-lZX}�'V��rtC��Nj�w�h~Y�wX��WG�%�����8g4���](M,bD��4-���8��"�t�U-���k�B��6���b�+��eYE�[�\pԈ$QbE�8�qK�3a��^�c#��S�(��T�q����r����Q@6Bƿm䴰��b~��i�j�PI5��fF�+W���������mÍ��0����L\Jb�D��%��������5������mᡶ*K�U�-� P?�@˗5R %P���3q�v5�N)ƫ��X��uM0;`OC��� H�Gez?:��B�%^Jeei|�*����=�&CB��q�@������U
��lT�r�����44O�ii��g�A���FGwD��겪��E�»�5DٵOTǲH���	��I���Ť$�Ɯ��gUm�����$�ĚM��p�](�1Nj۩v��MY+Z(���������b�iR>y�gȂ5�N(���}_���衕�S�1�8|�gdIg���7�G�"�J�WC�-k���I�=��i	7�t���� G�r�D�@LyT3�)�Z��$o�B��]����s��Os��x|��3���bՍ����G��:�Ȳ�e��N�N��Ɠ�T3O\��f��+
Cu裭�Yq�E�|Pq��f0R�c>�EX7�UH�4P���ǂ�_h{=oa}�<Z�'=�A��'�Z�	�=����O�I%h��)��0� LR3	�Eȁ_��"M������Wʧ�b��� I�sRh�ې���>�oI��T�.o]��s�Ȥ5/���H9��hI�8�^�s�ť������4	������lX6�C�^�W�,���RiزrM���~G��u�����_�拏n)�uI6-?f���Ѳ"��`)���%��h[rƝ��N�NIP_k���n@Y��N��ɕ�̛rNb-!A�/���F��꟮]��>_��N��u��}���[nt��.ٟ�[`�\:���n�1����1����iZ<���h˒���[s[�~Խ�Wv,݅ �k�\L��W)8W�s%���h��:��B��n�T	K�^$�p�t'��ќk��t�>�^�BM��j�mW�\[�j�� �F��Wuׯ��cK~"���L��e�.��K�
�s�5���u�N��m�(o�:H=�t13�:w�P]:�}��Xcu�n����~.��H�6�R6g�FG�2$�α4�2�o�@��M��+#�rFbip�u�C�ab-��%���u�iWd�-�v��ߔ)�C
a�D��+S&��䫞\���YG:���M�z�՜ +HMk^	��	~��b�;�kK�%2Qt<j��"�!�"*�I kt��O�T���v(�5��K�o�D����*��g�J
#��T��8���8Qm���x�	7
�%?+�V:L>�A���]��e$>Z�l"!$%+"1��9��pF�p8x�W�$���R�kBE`5�.�e�p��4ˠB[�����.9�n��%��#9���6��,��>M٤]����a"_��c's�W�:����Ӎ�]�@�==��hئ���"�pT��}�~��\����C2��f� {��lͫrQ
a�j�Em�m�`�N�n� R���T>f �8�cl�(�`�'fyVI����f���录7��d$�}�僖[9צ[��������۶l�� �:��h�_7��Q��8�Fl�i��ʝ9�M�?')ڎ�&�3Op���4�65�n;gl�1��A�N��}�1V�B9�ݼ䀮��(!Шϻ)y2TRy�����cS*��H*�`b���W�Q�"�2�Q$�`���N9�%I�6ʹ�6�<a�JOH�o���L��L<籵3���K���_sȶ�A��h->��QT�"c�ʯJ�R�� [q���C�3q]���[�3Úp �E��3��3���b������X!d��e���8�U���L�8�Ak��):Rq5�F���@ъŲ7�[mCqk�����D�=? [qN�>�&��v^l�,E�գ�7n�� F'C�y���r���3���c�M��s@R�� �\kll�9����FR�h��
�|�s6
���vA7�A�'�C�2R��ي�W7�ɽ��^k�e���|�����V��Vj7�
�����*R��k"�݄��Қ�zZ���(�<j���+GMsJ)�W���Ag�hcncӈ&.��w��:��8v���k���R(7�O��9j�	������nB��x���ڹ���b�������<���l��bH��Xw{����:A���Y����ӛz&�`
�N7V2ܣ��O�|�Ūҽd�ǏÞ���(� 8E8)�e�A?o#�Ķ\�5�e��8� �m�A^;I1��\WC�~�� (���*<M����o��'�M��i|��'/|��'?��s���.���3�u�Ҧ��t}��U|�@�)8�f9�M)`3�,`$e���ԦC����tk�@[�6�u�h����t��,�F���)U�=!�F�Ç��Ldz3Evҍ�f��f�-=�%8��c�p���!5R ���ҡ��	@�X�Z�|L��]g+���um=	���8fY�F�o����X�ת�$���P�����u�EB1U�Z:ƪ�i�ᶍ[��g�P	�ΐ.B�Grb&� ;������/��`YWK9E �b�E,�}_�g��7�jR:I��=�)�{��(t�$u-��ץ�򚡩|��r4.�.7W����ͭ�q�}�ś|&uQ.�z���u��eN���9T���ZZ8�M*"�0M�ױW(��ז�L��rԫv�=dD�oTDY��V爈��{�Z���}�k3eepF�0�B�̒B�"�0a�zHLx�h]	F��bd��bY��9h��k<ʡ+&p��mW`���ť��hG[���m>�P^��gi+Q����ʊ�I�Tfl%TJ>Z m�C�����$�V2S
���Im qx�R_8'�g���o�kb`*�8[���f��Dd"��#������Sf����l���q}Mr�9`z���Bb�׏�fB�Ω[pdw�N�41��Q�b�.�_2�����C��]99�=�01I:p�`��+o��8�у*e�Y��8�12x �fDYb�;IS�P����F�t�}�jZ�t>.��o+WM���FM:O�H���21M=�q
0ɒ">	+�DһCyʠ9���m]p��GR�W�2r|��+_q�-t��k5��'u��󀘸ݐ?.s�E���3~�l}�/��A���
'�!�jEX�p��+q�di��Yژl��B+�*'wh�٥��Ǳ�|�'Э۷��\����w���i�M��&cj�����A�����ӭ��\)���9p�T���?N�v��7���I;�D��tL���T��6�3o?�p����PT/\�(����� ���� R�(,�b<�k� ������XM ���k�R�w�ʬ�eA���'S�:d =\b�i\f1��c
/R=�Т;�X7�6��/�[%Ϡ­q�!��4:��(��"h��d��W����Ue4!ht�����	�؈m]{0ĐEG^���Y�]�F�H��_�e�����~۾���9T�$��8a9�n'�^�/�1���� W�&¹�FN@	� j���pV!s��d�S;ß��\�`��������Ӗ�n�:�₋4�N��}>�heۡC�H8=������'��,�=Q�
Yn�� ��=s������E�t��K6(E�"�����sg�qps��\p��� *���Z1�#�*ԇb�W�sw�?:eQm���LG���kx�̫\P�����7��H2P�m[+9�JJa��sWh�[�'=�����8d�7D��{�x|��7��vmӾ4���^H�|hPki�D�LMFR���Zy���������~�}�l^��\z�V���\��O�:4,�4�n����@�P�1{y���`=���7� � ����[�es����OK_�)�UE{����H�^���3�>զ���2�5�AI��M oVj+S���ܺ��8<��-k�kƨKL~��g�'��h�#�ܨu��e��'�ߺ^T�%<d.5��	��8s��Wa���c"_S��je���;�:�B��%�P��L>3�'W��%X�=j�cQ-��6�6a�v-�M��¶��N���q)�ÿ�T�dҧ���
��ӭR`Ym�xx*������u�,^������\qgT��`1n<�J��{Fx�bP�Smb_ё\QbE �#���j�!����v@�|��e�*�&]�qn��X��2Gb5f����%(E�f�!�^�H`�����EH<�����3�.4�2c�@맰�TEI��@�*?p�&)uu���f��4V�H/`0�'$�s2�k�6��+�����GL -�����F���
�e�kia�+�&���s�Zӏ��q�rN�}��y󫟻�,ݱ]ŜM�)3�)��O0gL�Y����7SAv�P�٧��(�sB�d9�˰�L�m�kA����u�>�s�@���XcG��r�{��^�����ކ}Yx�Z��F�v���h�cl�c�{��^�f��e�sf0��9��`1����\�,��7�l�jуB��̓�����]+gW1��Zf�c�B�C}�Ʈ��� � P-����5 �J�\��s��kG��:L��XQɂM��Mdb5��"��UU{]l�i��|��5��q�u���!=����izVn�)_�2�N�nμ4��}���.�����`�V;a�{R���	~	��i���9�l����� ���b��8���\��C��!eFA�(��sR}ZŽzt��e����L#�][����Q�A�K��Ǳ\�����k��{��2���3��z��VB�����JL��8�%~PҔ��n��"6�Q�7g����b��4���j���j�|�u�����O�85+Lz~�ca���9�a3��$ce�8��he[�P�
6�Q��6~25� H��#L��2%�Ji�8O-���Z�/�of����"�(�X�����09BX`�ԙ��P ��(�Il����:	���h2B�p�שH����{gK����C�v���UyH�cy����i����uw�Y:�F��~��N~C�K4j߮MR���� �F�i{}�������ό�1���Ee,�z�S�s&��_}��h�}3��@��N
��!�/X]M������T������NS�F)���ʵ���n��v���BÎ����Ш��k>?��Hw�"��:�@�*��f�Uhr��T>����e�L��j�/��FG�N�Ԁs\I!q!�\�Ua�,�S���`�x�BcfՋB�Ģ�e`$��$h3������3cyǸyf�7��BWf���򄰿���腅'���kM�Ȱ)�%�C�V������ܦ,���<v�`���L�Fi�عS�˴��ǫ'�˳�L��d�H�)��̓=�]&0&�-�|j���0���|6r�t��"+.�X#��+�U�j��r��^#_�F�y�ܬ�)2u/r��Z(W�t�a)uV7ux��%��:�$�Yri$\X�dj0{E����Qt'����C��-�n'���(�4N����%���\vJ����{�v�c�^�V��;��C�0yY̑�rmrg�`"�%�c�ޅн�jH4M�l(�5�F�\��튬��������E赬�jL�gQX)��G�!e��M�R IF���W��>�#�ъ:��lc	��\A����n�1}��9���#��j�(����� H���-�n;<�gh�P�H�I���Q��vZ��.*�p:x�oKst�z)v������j(s�e���Nc�Y��R�B� ����  ƃ��FcOP�<T�h���10}D2+���Q�)��,y�!�ia�X��U�.C�����lN�p8 Q�`�п���c�(�/��ʡ|�dC��+�?d�������*������̷?U��N�R��i�A\�<2����c�I�x
�����	p�z-��q<�B�#k̀�&���j4�'�Ձ1���64��N���l��o)�h�4ݰ�#Qr��%c3�?�HV?���N��d���rV�}�yމ��Łw�xx��.(�!�� ��%D���V�s*'�b���|���}m�������f�M>�J�H�y9K�1�&?^)���
�d��^,��&��kgpjm��+ab���u�����OR��$r�m��Q�*�@��;���L���=��o�~DM����>N�λ�c(�j��L��7��c�p��17Ѝ���Vx���t�pX�d)uf���ukC�@���X�#�ЄF3���11�ݥ����׬%��nbۊݬ|,ܙ��r�0M��a�cL\��y�|�-�͕���={�2L�J��ȪE�d���"��U^T��&fVPC�R(�;1i%��vR*�����Gf"�~]���B:� s:�+�^��jr��	�x9����qH*�q���흗6��8�ᷥ	�wF0݃�����?H�m�.�ﰍ&)�,~DX~{~��n��e��F���K�{f��y��8q����k'Ln޺���������x�0�@w��M➷��A0)�����酄@����9u�#Rv������X({l�-������I]$�ǜvp@��s�#_�����[	A`�\�kc�P�?������e/�y�����r�l��RzXe�JԔ>I:(�`�����>��آ�bgO��@E�ۺ1��+�gC	����;;�n�=E :F���1\��d�vd�����`�Ā�8g���:J���&-5���q�Q�4?m�p�
jYS,麖���reꀛC�Ћ|Գ�_�Z�g4�-9��7�/���)���qk//Ō��GN-���G��������u�p0rP��דkk2��2��#��P�e��k�w(�GK��
>��Ep�֭[���c���7� �r�j�~��,;��\D&N;�P�)/�����;����L����ĉ5����1Ž����E����U�WX�#LD	�P�zN蝢�/c��J�*�����B���0PF2��<yq���9t�Psǂ��db��)v��Y|A�
�#�9�D�����'/yu/�����ǜR��'���K��Z^����W��Rx������s��?$���!�J���pj���쯘�֓2)z�$f��]˨�=m�>�1�4��%B �ñ��C+�FvPa��٪eYV�=w��&�z�"����hi�p$e��V#��DK+�����+�*�όD�DPfpjI2�W�	�(.�����\>�4�s�G��*M�K;R��ܗ0����_�`�G���n!��(�BϬ�v7>I����V��V��/�x����=�����I��:��R��)c�6}�7tO\Aq��N�����<.K�v��K���7L3��
5J��A��n.��b�\q�V��2m���a�� �L�#ٱS��ŖSs��\i�~�نȗZ�pfk���n����[s�*��t������b�q�D�0�Q[����@�,�Y,U��0�D|��M��B��2�PMO֠e��T����/�L1��B�wD�[FJN�őu�H���1&���œ'Oܻ�@��CA��qX5�>6
�1�ґ/�ڎA�"�=��_�u�?�"u�E�.y�	 C�H۱GÝN�M�u�g/6}��R�5�LSO>�$l�e�'җ�&��'��6^�w�rm)��I�	��ݷr�0���>4(�FƠ9/X��z-e�F^˸W��M�����(�����.
��'ǁ�X�S�X7��ᰢ>�˃�s��@B��H�� fS�C.t��)� %&����C��_��C�C'�#�7@��Zeaܿ3�wT��3�GQ�'Ë��J�!mU����W�!��Ԏ����RY�'����j�.���5���U��h����s��5�$^q��r�iMQ�n�"�ţ��α���r(Pb��fC����NÌ���E?�Z�(�%1m�G��J��q9�������Dd?"���W���voi%L�#6���)j(B�v27)(jF�r�r�`�Tk��L��8�B�iꋽ�9�j'��F�K`b݃J��ͥ�*�%1G٨Jt]-��^?��"��ڵ񘦦���Â��$��W�/x��w:'���7�=5��A?�24Y!��0��I:���:���6y:���)]XW^�*eق��0K�E.f0s!`�НYQb��V��tv (v����/n^�)�'�DЖ!�^���T�Bab�׎�8{<�jkZL鿘��JQa�SΎ���ov��*qhF�b���C�4}z8�� ���
޴4>)H�!"&��&seH��`�xJM��l㋺4�iㅁ�߰\��PQ���Xu�1*h���iF�5H������[���m��D���'6�>3��:��pk����dv5��N[ϛm+2�ZZg2ڳ,~s�I���
�l�q8��W�d<Io)!���,��*�
Z�P��0V�O<��PJ׽$qi�ʚ>����b��cx�˲��(T14�`ǿ����������GM�b�@�ٿ���C���x��l�D�^���>��=��V3GK��b*ǲwѓykN�F�L�Vn�b��B}F�Z��d�);�_eʵNA�n{��^=#�+��Z_�u��x��9Zb����|: ,���u���P#��fL��#G��J��)�0��׉�	�4�[����LN$Prl����a4k�2
��cb&˘ԧ�����Ӡ��[V��+qeta��L?���>���#%qj��E[�g�5��H):��i̦��%��g���I��)v�.ү�[_J_~���rl��۔�<�&QB@8�mN���u��G�EȤ^�0�k�sS?�0*J�3ue��w���W~<Q�u��e0�4}���L6����L�I"���"Q�j�$h�P
��o�e� �\R��41�,l�����/�LL�K�T|e�ZyE��0+�a>?J1��_'ԣ�a�D�Q3�O��ob�$F�$��i�J&�gZ��:�E���g$�OS�P�Dbk{�:�qu���X�̜h��+kQ���o�Ηr,.X�Ǝ���f�Ʌ�a�0Phڨ�^y��)�d�h��s��wVw�;�(NL�rY��3�i701I�#�8ȧ�2���~� e�oA��ï1�.{���zEm�+W���Yб��ǛO�D^kk&
-p��^R2��S��Ŵm�0r[��`� �����l�E9��k��g<�b�t��Nկ
����e�x(4��>��;�Sa����I?Ōg#�7���F��Uc}��O�񛦛�[F~��Eu���7��X�X�Ρ#s5S�؈��E�8q���ӧ���=L����+T9�nO�v���Ż�q{P�����n:x�[T:������y��2��p��ڼ� �g:-Z�4񥛑�eٯ��B�����46a�M$y���9K���y�ᢺ����ʂu2�i�n�yj����1P�E�-�+ˡݢ^�j�Z:��&�%R�;�+�|ʉW�kG�߄�v��sZ��Yx�	���r��ջ@��/�O_�6o{���kZ�f#K�qVp*������|��O�F*����\;y�.Ӧn�}e�$� ��#ŃJZŐ7Z���y�+�k*xR�.*-�����x%�6A��mtLڴ�8H�(}���~��R�@��ENw��S;��-Q}Y�g<qb*����RP�
H(*:���jr���3d��y�i�����������?�h���f'���!®̤0�Rcb�ّ�ȉ֠�-.�	,��>ɋ��n�2�k����h�h�E�]�I���4ࣘ���:��~�?C��cZ;�e,y%j*����3u����@D& B��L,�����WŻ;{[����4�!��Y{'?��5�����!�F��(OLn�u3�0�߸ G%�^�X�4^�#���j^yc�̈�,��,`b��g��I�H�$@�t,"�n1wtzG�JI�t�j���@"ɯ��~���iw��&�hQ(h�8�6�;�vLi)s����1���@��k�d_ϘN�7:
*�/U���Z\LV\Ӷ"���o�P(E�:Rt\���B��Ԡ��ݸ�o]f�X;��iwaV$17(���eQP?vW=9��mհK0J8��1���U�x&�� a�"ub\�ts^{��N�փ#�.Ι;z�Sv����T�5����2Rz9�٥Ce�e��Bێ�cP����9�I:��p�ož�Ȅ�[���l8>�cM�)F�bd0����{�M|m��p�p߮m�p�4��4�ۤ�CL���E�j3e���h��?Q#�����g$)F��Ć�����<�/͓�]�	=�Lh�1�Ŝ)i9���z	B��W��<����6���Ӿ����I̬m'�=^�w�D-,vJ�7��y�����a�t��dk��Y�
��]�3�� #"P���m�)^��z#b�*:�_���C��C}���]!�X���b��e29k��=�Mz6�-��Bg��<N�WyHB0/��π������&�H+��1n�>,R��Ί�Pp����Y�˷|<���`*@����N�q��Jl_�2�Kۓ��1�|�)%Y21rK8�F���۪1g%
9K#��	�n2q��RC�Ź"6g �T2$�%��}ld�CLf��$�_4�*�j�aT�T>�zŀ�mX&��zL~oʃ�� ֨K�0�$l�z�iCJ����2���y����R9>~��J��=�sp9�qg�ё<�\%��CC� � ������L���W2���y�����L-c��S��9�G�%�7��o1)��N��+@�)��N���7d�\�uެI�rB�-喬�H�/��:ڤL���C˧�!�ߗK'5�5_��ehx���kf<m��"�_+�=k|L]�?E�� ��CLq
��.��GlǺ�Υ�F	��i#�q_n3&��k�>]���'��K�a\q��E]�&���Vc������hm29��AЎ��f���K<�¬~�5fv�mm?1qi���3�,�4m��59�,f�D-�e�6�kF�|�蚷i������%�����^[: �Ĥm��	F"�b$���j�O�� �����@&Gj$��,�����+�p�xm_��x��19���h� ��޾)�P�B\�$�$����<���>_��$o��[��Ve.9��׬Դ��Ƿ������N��X��q$��IᕝU1N+�w��VU��H�>�dVȒ�l]��oCz�k6~;���]19��[���j#�Hb�dH)�� ���ށbZ�ȱO��@R��c���m�n[J;?���do=�6S�/)h��j��s����Q,�� ,�|^�؍c�CL؍Cu�_�P�BEf��8\<cևq�+-�-�'�m[
GW�ӈ�����B1%;��Η� ^6_��}�=�u�j�M�)EX���ϫpŭ�+nS���ͧ&Wӏ�_��@��z`"=��"`۶��g7�� B���+nbZ��&���U�FMSí�sH��[|&�3Q�n��@�^=pJz��ӝ�pC(�<i�a���
���	0�L>||����! ��E�P�(�9:��-SL�it6m�/�K�צ��7W�h`8vIή�Z�`����.����"�����E������0�D��!6O7w�+Ki�<�nA(n�k)N��b����I���OH�Q-Ot��=,Ԝ����U�H���7\јX�H�7Un���������_[Y�B3�ձn�|�>�X G�؍��f,ma���>�K�6����nz�١X�m��ԌN1f�{������K��ڢ��CA�|�^�q��WrF�ѰCu��֧vrI��m�&%qJe�/����{���x�^��]�5���!�~bp�	�q��2���_}`b�9#���}����*	*'.�8������uB�
n�:e�zʖ��S�4�l��%�ʅ���Ln�+͗�R�p���aJ��8�8�ֆ�A�\8L�����M;,���M�:8�3H�o��X: �#��Y��m�6o_�O}}-��ݽ��=�KLE� �PͷC��1�f��]ݺ۳��W�����.>)�	R^@>�CƵ�ֿ7��6���A<R&aU(Ȯ����!L
5P'}.qA,�g���TOLm<8��E��T`��;C=5�&jԡ$�Lb⑜m��Ԋ�6%�"{c���p��	����
 g����e����B��m!��Y g����>'cm��\J<jO�����b���o��6�������6�E�Z6#ɀ^���;�5�H����0E�����pµ-fmW�{���(�3Y� r�<����"B~@�Yi�,��BōЇ�hњ���?��ڽ2�<	�EK�F��ge�S$�h�y���C�������+�&m#�ɺg�ӻ~}�<�,�p��Rx&��9O�ڽ�fH}��@m���b路*�\��3���d}ᵞ�$�eV�(2�&(B{�`���8�D�D�����9HU��h�V>��9V�a	�1ءV�f ���X_UL�����=�W	��i���"PP�ɗV�KB���� 3@̿ ��7�Γ��pL�Z�X�"°�=\�e+���5t���o���xfz����Zd�~��ն��k������s�w9��-9�9]@���P�$e��1��fԧ>�S���j����
��
NY�r��_������f���_?1�2��b�a�񼚯2�4��5O��譵jb���qzQ'���u�:@(������8"ۼ� C4�A��d���;'b �� �5S��߽xݞ H]�aK��B֞�Y�nkK���5����v)���7�?�!�zc��!Ӆ1�+?���K�.�w�*�_	�V�#�:����ٯI�-f'�k�UQ��va,���ӫG�~��]Zb�^�����6~<�cf��ǁ���EnO_c4\�DoW+� ;��yW-��%���'���3�=�w��OV*�|
�f<c�56�Pt,�G��~[�z����!�k���*y�-/�
��T<�၆	soJ��2����v@�  @ IDAT���RcH� �48*�N�/6��'���+�	��q��w�tzY0�0����W {��jZp�a�xʎ]� �^Ll��kd�g�x ��ˑ����� �����v�����7ϴ�K��IE��'���8L�OS�Aڴ���:=-@mp�Q�m�	-�1|�A�f$ܲ�ȧ7{5�@�pcc�+�����6�H�@��L^���d���������}5��(�j�w(P��?���&���
r 8��R/�p��&)&��i���x}��毄6[�t���?�ρs����\xC�b�7�#��.q�t�+_�������k��i=-��ז�;-I��+����m��O��I��WPd�h�1t.��Oo=��2�9Ƅ��}mk��\_�����<ܽ>� ^�D�� �z`S���M��=�t3D�պ�e�w>�/:vb�j
2�a���S��/o�F.%=C��,�҆�9���XL�
Z�T��y#�u{i���|��^���>����Эnӧ(�L�o�h}/k�H@���۾�5�S��Lo�:�w�i�&H|J�: h�Hz%#
%�ș���f;;/\���};A^.��mD���+�ap�]�U/]�*�J{E�Z{�5��MK�!���B�~B�U	V����i���{������@�7mG�/��~<%h�q�GS�Lh���'2��MzQ�,� f�"�ߎ�->j�,���Q�y��b�%R���.�g�,=�ԑ��@�$�Oc��ʿ�}�C&���&I�8���.Ý��g����zF���;�S��9*��*@K��>|�@�1���r�۽�O�p]�_�ڃ�&Y�n�Myp!=Ob
ɔ$�0z�Q^���m��n�6}Э�k�;��o�#���L�V3���*�/]�,�;�k�W��[9���HMƱ`���k��1��ʌ�=;i�`�=��j��YG#1�3��dF�3���e@��T@t/ߙ��e�L���A �G�Ѷ�T����|���8DG�ǈc��!k1A\m�r��{bz*����1q8��^����_����sTSm19mm?��W�Ǒx��٫W�
�]�����/_؜��r'.�>8���mv�B�Wk�CC�c �eo��q{j�T��j��߲��J50��'�T�T�>�b#���Q�j��釢���Z����,m�%9#�E1�N��Ts�4n0�$�q�����|�����ׁ�5�/�0���v���w�T6>��qo/����5o�x��}Q}�i��@���U8�5^�+��34��V*�i���?��R�#��9rU��n���T��b���&{��7�W&[�~-R��\I���ܨ�ݶy�p�w4܉�vk�Ss���j�ڼCr��0%<���7|{� ���〸�rO]=��O�u�&-X1�]F8H������#���J(�9v�S��V
�% i��u���3d�D�V����̴�a�������.�&h���ߦ�'L��+,�1��jq�ԙ���c���2���ՕGO��zC�c�vbU:F4������r�i<<���㍿j'�Ȯ�t|c��-#:�b����㚞)���Z2xk�ߘ�9�@yIbL����铇bS�z�k�X`(}3�bbO����ٷ$��$.�ϟ�%�\H*�l�����-V�Ўwc]޿5���B?k����M|l���^*Y=����S ��g&ԌsZyV�A�6�5ml�m��(��mQ��y�@Ky	%�
�u
�]Y����4mq2&�փv�٦ڽ�Z��kX�Y��N�fn��D�OJ0y��G����?���W����^�Z����u�d<���eg�=�Tg����Ƴ�y�c���ޙ�a9^Ɯ1-�6<L��` ��Әa?�)�1K���K˗��)Zjd	L&�����1&^L�Ӗ���=��߂�'��oF�ڥ��x������S�t!���e��r*P��k�x݃����{C��������K/J�L��8��#�G��P���3ڊi�gtP$�+c����G~��xr�����Կ����u+�k����}�=�fh������wq�o���dx�A�Ҫ�IM?��8��c�,PJ�1����i��j�Ú@	�O��ԉ[��q�q	�3�Ӭ@2A�E3��'O����=s����~��gΜ�4��x��X��g�^�p��]�xb������g��/�����]y�ki��y1ܼ�i۵���W�~G����W�q�MK?mܘ�Dإ��t�Ґ4K�o�ի	4�e�k9��mJ��iO�?�\�lh�]�3��
����?��������3�._&�/]�p�I^��6n�	�����C�����Cw� ��s��{a��u�#e���'z�H���V�%áW�O�]�ѧ$��DBC���~iwv�A1�?}���Ryũ�5	���[}�m�����5}���?=�-���[�!��gc�Y�p�Z8O�6���=\�E�Oof�����ڑ�й�ׄ��q&0%��oM�*}|����~�!��uz���>9u
}�ٳg����7~�?����~��޿��Bu]��v2��k8}z]/�NI�9v������WC�-#X���C@'�$����Uq�_����T���%����G|{� �y/ۇ��i��	���B�6�H�m?�|�}AL��~��2^��V���I_��J���C|z:S������/����$�n�E\�z�NBE!��R'~�~���c+n�j�f3��y�X�6*J����^QH2XHs�N$7�sT{.Fq�F�s|llӭ����4:P�/����}zh�Y�&��i�qW�m�L�,q(��K)*1i;�4��W3�����PF:�:
g[`\��b�������л8�
�b}S��G����q������ӏ>2:T����o/�a���-����A�:C�Z���]M1,��U��|��n?UO��7���r�/��2L;����P)O�[�O')(͘[؃��Z8�s���?��׎������|L�R�򱤧O��p�҃{w�Իqm��y�kcc���s2���C6�"�pU��0P�ߟ
��i�������s-v6{~5~�j��V�6,���C.;�@m�FSa���>��#w��	�M{zg�
�f�1`�a�<�Cu�UW����R�qR��it������VF3��<c��x=�z('L{�n$�/M��XB/*�PY�[<�5^-�i��4�s��^PPW�^�LC�͆5�����8Lj|��G}���C��y�ѣ��?{������}Ԕw�Z	���6�#F�˶�tV�o�[t�5��m���Pz��>|������Є�p��2�^��D���,0Uݯ1�Q�$���(&7���@���+
>�45rF D�˗n$
�Cxt�hШ�C�Cp���Q�"K�(v�1�{��Y/�"���_�~�tl���}cV���\|\%�w�я~������L?x���x��,&��on�'/ٳ�"�,W���}lp���k�%�4edK��k���638�ө����!N����̅���"�x&��f�q�ʐ��g�Xs�Z�������� M{�^�I�ΩA��An��s���Aa�:bb7ݫ��#<��C�2��iW��~M�j$���9}&Ζ�\�Ue��8[}o������~s�扵�ܸ@��6���)n��W�#�c��%��鏠R��ǃ^�H��'6v�v�7a�kk�!t��&v�Y'��a��y����Ʒ�5�D��a]p��j�)�=�:�RCy�_pM��{� 4��&��4E+)j�0uI��M�=�!G�J����3��-ڨ�>^��Fw|�Ȍ�l^*XU!8#�觾�G�Lx_8����n\�[�����_�7�9{�����?��J��V�?$]�C+[m1YB��P0:�B�q9`F��rU�& ���R¨�'��1�負�E
!�c���u�����m�o����#��8�v}N��5VnO����4m@�J�j���27U7��<����qa�	#T�h��qi�\�����F� A=�f�xKo�;�+]���ބɮ���}o � 	�wR\�M�͒�pHr�5��D��{��xb��x~/�Fϣ�Ѷ$�"�q	� �������v��yN�<w龽�z��v������ee�G��bzY�K�b��92��<�m��>�>w�_����f�sZ��`�R�3woai����N�t�J�
��g��pL�����{������4����$�����L�qa=y����ke�|��~�Z��u��m�W��.D^)�)QNX�B9��l5�g�},*;�]^��txg�:���T��vD�]�U_����
-�PUg��@��	����1�[�z��4ES��]���Ry���m;c:W"n/�D
�zb/�g�ݸu��=yJP�d��	�ޠ�/Wy��ݰ�gtlx���#�<r��5�L7>Rǈ��s��?`��^�(!�q���&�>jv�J�t	��`��:�*�G�ʶJf��_[�Q"���?<828���{���
s]��5��ط�&fe�h2����r�
O�ҲY�TOH_���}Ek�{�[wj�|���߾����}���G!R�,��YӀ���k�͙9�0��$�*a�Ǣ.�|��'O�����dZ�`��M�3�'�*�uk�h���ЯL�X����
�8��4�G�
�����h��z�X�?���q���.�߼{70��V_�%J����8��ro�Yw-�4�?��G2�!#J|"|vw�EQ��o��������L�^y��) ��"t���?��7���8A��`sn�.݄#k�귩�\��פ� �I��o$�	|C�7M��w��� �Yɫ�7����mT6��h�U%*���cG��]�^�}��n�.H�\�������$�޳n#�,<t�a~�硥! �T@�3��6��d�K�O�I����ȯ
0��������FBZ�ܕ�XkW_^{ ����̋|g��[�̐��y��l\�U|�;��y��rp��Q\�� �����ȿ�������~��ə���c�8.ٹ�TleҞ��a������Y�����d�����G����I Trũ��ɠ��vd��G���&+\�H|G�O��
�K9}�̩�z-��`�	.����S�O���r ؂��F�9pf͕7������2���>�CƂSmN05��%M�<�}�=D�b��P>��]�ll#{T���I�C�_ �V��G�o���������c�RД�m�·��u�� ���;w�0�㞁奥���n\F|O��Ǟe��A9�m[S�\s�;�68A���"y�9�8Z�2|\����@�L*��:�ݐV�on..���W˫+��H1�E��H�W��}���$@+��Ѧ��`H�n##�G�rZ�6A��&�1gJN"ّ�擀�v7Ы�ʹb��M]L�J`�C,��<��m�7�w6�jo\�z��-�����p�,�m�`���=��^^�֙=}��AJQ�<N�rdb���3���"�aEQ򸸛]A}����T�0+�guQy�� j�haH����ͭ,-��  �d6��t���\sQ��%��Y8h��V��NQλ�V{���2&0�����ʈ�3?�dlh���x�2Oԅ����js�4E�k-��X�� �O���]��/!�\���y��ŵ����\7�ap��kk�����ť�s�oaa~an��8�����H�d�q`���뮜(}�
�k�f��xySW��h�65����beAh���+ҴI3 �R��m�㡄�*.2���T!l�6f����`4:��(��8'�Ǳ�2> ���$U�1|�'!<��; � �.����)��.��� �~x
vy�Ǌ�����+�-\�5#>0P]ݔ1hR~�V�z�i�1�Z��m,<G��Fk`��&�|َ��	O�V<H�D=z��x%%�!M�[���n���I�U�a�:v2�oI&LӘ�Ǫ�Cut�*�#�.�د3���o�y�K�/S<j��V}k���	�3����>H#����� m����hD�������HS(SH��Z���D�4�Y����Z��*e�y5��v�
�
��̉��U:^2�em�������@A�0�-e��X �<���L�%�Dᗺdف-��c� ;�r����u��zM�4Aq�s ����4���\8^)jG����GMH��m3�w�����I}rZM��8�<�_O"~�\Ɋ�z�JO'�m��3�������<;�nQF�c�g�[����z�һ������]@�s�\sX:�4Ĭ����!}�r�̵�C��U�`H���c#���R!G�Y�l6חu��5���j~�u���=qb�5��5���Q��<�&}�.�սx������=X��#a��o�Ѡ�4���ࠟVp�d�X�Tc2+ɌsȴXU����n�ee� ��+n���xφ� o�	��X���*�"0��� ]Z����7�}�N���%T(/cW��/��d#(��f#�V����A�������A��6���S�N1ǖ�ᡮW?fv��W>����������L�kG�OC���8�Se�c���<<ҷ��
�_�`C�qw��0�@��.�iN�E�m�HO ,vD̯.M_?%d�{me�B�	��
���jZ�,�R0��xe�򾝍Fa64�$}���8��H�΄_�K���	R����h#�lӃ�	63�yu8H(�Jv�> a|�,2��i�QI%>E�i2�H��b���-(�9e��A9. ��'"�`aK����R�q��(�;��<.O�{8ᅦ�ɓ/��=�p����ׯ�ϟ���<7w5�uEHb�	3 �Rrt2R������陓LhLMM��ii��������w?��5�,Z[k޿��YkC��������벆2�<t�k�WT������u)?:}��k�=ͭz<"0��=��8oj��<���_ į?�'�W[�Iԓ�3M?:�#��Q���A9ǂ N��(�`DA����1*� |�l��l�5�>��d,�3F#]B]/
���6q�DtyP�k���(����xm��J�?FI�{�#*#�b�cD��ˀ��zs���C�=������[�n����żB�\��8��E%�g�8۸	rHv�ɕ���e����[T*���
�Ӕ�L��к��!>j�c���ŦÙ$���-��T�:t�M��B}���P�'2����P��%I�/8H�C�O8�zb�
�}]C� $�dr,����"�uz��%0p���,A����C:�xi��[����''V���O�����t��K ��p7��1S[�cjm��ݕ�Uo����/�ȍ���3zIn��j0϶���ְq���v��F�$#��}5��N|UU,�J��I���-5��%�c�@iջe� ��I�����8#JG�+Zr"�y~Ut:�*b-�j����T��ؓ2��>nȸ�f-��_��o�P7k�i戮I��f��/�EM>�¬	J��>��]�A�=��~��G#֞��Xv��{w�D�Y����Z%�7��@EBw��0Y���ZZ^��d�2�!lY"��bJ=��ts�ZJ�]��Ef0*����U�� ���_w�Y��{��X��t<��J߉YƮ��2		��X���܆�t�p���$2V�?�gw�z�+�u�S�O���d3=���Exj�ڠ�L�T��CgϽ��kgϞ;���Xb�2���s<1u�̙���U6��\��7�E�R�nc��cZ�{@�����֚f��
����%�V��k1�cƩ M�[���V1TV��	�eJj�����uF�j<�ֲ�I���&��5�]HA���,�^���Ǣ=X�jN��P���Oa�V��v_��Ve�rxi�av�zyر��p#�pJ(x��UԊW/�|,^���'��F�51F
w����$�tk#�5�"���`��Ȋ�<������l�]1d���@���$���qB�!��'��xukՕGt0�-���_e����Y5 ���P	s�գo�߱RD�B�:�)�Z���qq��YK��߼ߟifB���]��\�N����������gwS�:���I%�}��'�z�g�y��gfN�~����9�U�ԘwgX5���ZB/<zᗿ�m�倥e���7�۷o���RS-,�*:�#�.x�H�O�Ō�;�,�� ��d�Jy�����W8���xW��]uM�%���k�]}�e}�8�Bݧ�{�n�0�F��������?�FMlb�s65y���n��}���1��~��v0��޺�^�ך�ĵ��n�b� f1G��G�k�G�F'�T!��s;���
�5o7K��U����3�	e�
1c ����*�����4�g�[Pv���aaʸ���~�����M��yz��6��;M�tn��L���*��;��Op,+��'S'��/3�a3N���+����9V�\Ԥr����ZŹͅ�ȺV��2�κ.L�A�C�D�g셸}d����v�.���ꩤ���_a�x��䈤S�U	w�ϓ�iE�\-l#$�]d�"hJ�3���n8�i!ꈅ�m#����i�d�6{0o@!���:�&��PD{ �SO=���cb��L��1p֭f3�½}����͞O?�T��:tw�����d��8�:$h4"`�BS������R��g�dZ��k�lZ��1ߪ�P�p�r}�槠��z�� ��V�����O7��Խ��΃,����pU>صZ�cEEcG�ЫqS�Z��Z4*n��&ƴ(���ub��&}�Μy��ǿ���-�<1���"�`f1g�;E��S5�啉9��_#F~3v�����]�÷����̺*�s|2�^�;y�9�+y[�����5������RT/ЧR�X��FDz0��^��Q 6�`��r-�a�������in�7w�b�����W����p.�2����Q؆$��%M�7c1i�Y�c�����.��>"��q5���$�vH����\w�U�v��!�+!g��,H%
w�����2bQD\^��� (����ư��j�	 "�Se&8���7��2��:�Ɨ�ΔC�Օ����{8?����y��H�;vC�-KO3׋I��<���XcO���h��pd���J>¨��ː��
p���b�n�wY��Ѫ�ۚ_Mt%Oy��"]gI���Ȧ/'�Pc�I���D0�T�r�{e��o����n[v2�����R�z��
��m�N6����>^^�LR6D�>�˵ݞ�K��&}B��1ёݤ���T�Ϝf~✍�(l����"���o[-*ɡ��ǟ|�Bmn6��[�n��mz���g��r����1>��n2�&��c_6�����6�K��!�X���-�5���F���Dgg��ݝ�+�W��������@%EV���6Z!Q�<՚���'�w�g��T+��A��B�b϶DAa��'�$0������M���-�:L��u�8V벭���w��Ʌ9���O?������Zc����S�����l}$�����*�V���$y~����`\X���p�Z�:�o��.���k����?l���b�?�(�FE�#s���~C0IV�X-v��eG[���mY
�+mb{�����` .��ۡ�L�a�}%�3;�e��{��T�>aN��Uŷ���S���?5{�4�>����>���g�gO޾u1�-�
�bO� ��¦F������1�Ͳ�%���|S;A��J��:NC���f������#	B<Ühd#I�Km�)}�Zo�
�Y�.h����g� ��e5�0M�R�V���&����髲�vq)��7�޽{���u�Ӟ�>��qY�"s����3 ��ܽ{O<���+���u�Qf��NVrG���A }+��N)�CW�lRE��Qv�7�����ۮ��ȧnW$ٖuߨ0^�����
���R�����<�?�6v��GHΟW�� �c,2W�}i��Rq�$h�9ش�-��ʴ�SN4l��F�l�!2�5_�s��ot��"���|�\^Yf��������>F�5��zG��u�E���9�<U	���+�P�O��x�x��(*5
pHuwz�R�1_(��+ fF��O����َ]O�s���6�<)w���m��R�2���]��+Evy,%���d��ב��������c�,ma3hzN��G�d����C������'��V����o2q���S(N����ϑ���-SO7Lrg=[�gΜ^\\ �^&_�����fLxiE��jF%S$U�F{��r�)���{/�\mq�J�ϑ��&ά|3�V��A�64�3W���GN2F�S�Pһ	�npM:�z�+� h8\�@��T�� ��$�w/�v$�<�?R�� ?Ԛ�d"��PL�@D9�t��!�yc>������_��׿��?��?y��+c�����J�U1��l
W}�5�gO��ߝ�`Ld��-�a����3�A��Xg��zTt��H�zm�+Z��+��<69��v��O�J�C�	�9/���BݖA�Ӻ|�u����K �0ʩU��=�9n�����h����N�P(��he� >P�>V�l���_^�m�<�a���h�+��0�Ŕ�_��_���!U;�������t-5 ��0�����Aj��Ȍ8�T���S�C+m�¸b���;tt�s�����VU�q>��Ҁo��-��2�>����n�}f����g��[��L�+�4� {\�p�[o�5�f��!��������}}g�9=9�
%I)L���W�eN1PF"���{~]��Up������PR�H�V(��~�R�%n3���+����rMA$�|��Y�FB����w���?�iFr���@���!��#�ζN����s��20bOe��_���_z%��m����pLU1�]�"^����lנ3�f�����ҿ�B�/�}�d�7K��ctM�cUKj�ȃ"Z,�c�@Ѻ&�'��,9�	!���鹍���fk.��Ϋ�w���W���2�|����l;gwC��:* ����Dl��Zwz�:]`�'�4e�l�� �a���!-1᪪ϟ��E�s;��k���&��x�lDi�����p0�Tc-�[�0X�"n���'~�x��^�V��5F:g�¹sg�y��lv��~����5=��|_�����m]����Z��ڵ�zB-Íp�Jw��`($Nc ��En|� AEU��p�_��^�����t���4h\�oݽK�ʂ%7�1�D*(�Q��>���!)��Q�6l@K�PRz��\B��	�lߖcڇ�g3���է�`���x����AO�0���d����.b�	[��7�F|P�b5Nj>�9���V�2	#2�Vu��(����9��иq��n������r���č.��q�������+���G��9Y�~S-�vK��Gŀc��L��[ͦ��F?
��˸:%S�k�O�՘lF�1�\bz%�p-������C���	�)�R��qn����~a��*���Ӌ��Z܎cr���P��o�#\�_�D(Э|�&7�#nɦ�nxZv��*�
Mzt�>�Kх]�A%e�3	s/7�\P��.}L���-H���Ro�Ք6��ww�4_���f�������~���_���ׯoq�����**��؂A^]�� O���9Q*z��%�>\�A�?d;:=0<��jZ�F��yqu�n�
�PBh8�O���CR~�r��;~ v�	�1� @����grd��D�^�fl�#����K�U+ڤ�)�Z�@�aZ�(�_���a�����e�G�( ���0dY�0�W��"�dG��^��;rE�`m��+l*}刧����|z1��<i��&�j�+�rY�_�p�,GB��V%�C"�{:*��Iډ@�{���������?�w�ײP�S��F"Ԝ����2�*��+��$֊7M���A����S'9yå1K�28�g'�� I��2���b�V��	��)ۘ�����M����}}��� e�D�oA�f�>}:��Ξfm� ��B���H �P!���Ow��Z���c*7��9е'*UJG@+n]�E��	�n� 8�#��]���RF=6>F���?�������t�-��l�t�-��C��p�ǉ�������+�k��5yԚ���z
��ۭ��r|\�U�� 2i��a[��I̺�m�#�"�G�%�dj�u�5�W�>u����-����ϩ�S��uyf����mF�Qa��`Y���?X}x�#�Z�P�L�8s@r�!�D���I������1(�ڲ2굂Y���LU��9���ۀ���F��+
�w�-��ŧ��<�!�J�vp��s9IH�b&1+ �1<t�£Th;�=}�cA���?f��G�.��׹	��J�ն�7h[2g��Gu�Y�c���P�ZBrU�\p�6�!�XD/���(F-�䥭U�3i� ����Le")Dc��z-Dæ;��F�\J� ��krE��Q�n+���
��]�έRc��b7��8���icu��Ȭ"Q�(2�E��@�S�y��APwxՂ��Q��N�u=V�v�l���x4`�U&�H�*D�ʑ����4J�}��N:!�J���d��x���}��'�/-{myk�R=��|��ũ z�k 6���.�w�mnM���@���'E@Q�͔R�}��Q}���N�Ɠ�Ѡx�<��j{�[�`{g�¬�jaZ���M�w���u�8m��2&iL�� ��QZЫ(6A�nƠ\4���>
�d}K�ę [̉Z�
��5�� �nJ�y����c��f<�ڮ�*���L�D®���۳q�8�^���G�$���c8�.�Yd۞��g���v��`fs��pa�0>5���[oڞ3(��m
LM�"F]�±�D�t�,��0P���j ў(��`
 �"�J^B���bF�0fyuء�|ކ�v�cA�yM욤��C�m	�r����OK܎���O��
8	�=�'��K������}�I�MH[�)��H�j�Aß"������ @a�`E`ULLL�"�կ~��mn阅������i�X8������X�V%�<4M���%������QN=y�b��*��h�.w���O k�a}��2����'�&a��0����%������ٮ�Y������\ƪv՛�d�K��ͼ����U�
�"���Ƨ@�#�a���������x�M6W0Q	��8�iU��|>��L�y�nt��STu<�S�ز݊�Y�0B� 	
7M@����
A�_,`�6kw=Tr��ߨ�zm����t�>9?ݘw���b纨|q��\�<C7�����İ�ŇQR��:b��٤7�x��^{�5v�OO�����X{:�c巿��;f����u�fO��1Ӝ� ��y> g�a�+Q��V6V��ě>��;���,���+���^����@�c�!0T�7;<�PXo0uz��	dA���ߚA�#���S5��d�;*���e�fΑ�Y%�"���x��ҋL�ʗ:L�_��UpA�!.�#�>j'��(c&�''�8��������l�E�L:=��-2�{5-��(SZ �e&��.-���>�BV�Y`�J�T�����.�(�;�����-T�_�2<,�ۙ���fq�[�/َ���c� ��Ov��Ii\%���S�~<���n� ��Y>���Av`�|'''Q���|����_��/|�W�sf�ʡp�I2��n/��k�d��f1��x_�/6�Q�]�����a��Nh���AG��$翖�)d����5��
�>���;�\YgW�ru+N0�U�#��P��,�]���~�ǸW��%�c��ǡR>����~��O>b�krjr}qEݓ�W��m������Mɴ&��>,��^�P�o� ��sj<-���ھ�ԇ���l#e�$�䟩��\��Z�x�,%V�N˒�6W�S�[�������NR�#�1�Ҽ���W���-�_lhg�Ps}��D��D��1�t�C/*�׫w��STs�Y��ۍ���'��<�-̒bBc��w�(�~:��0d�^&�@���R�Jx0�'���V�)�(BZd���	�?���Aq�vBX}�����<�575��u��ZKg�>I8�Ob�b6�FJD�d����W�����k7�^���j�t�}�#W���$"�]G�c��g�}vc����ϟ���!�9��[{O����<g���I��1�wq㹭=1Eِ���l�8��ߌ���4*��'�<?�窆���&�ϥ�yh��ңtfrL�ќD�f�����Ju�t
X�2&��̍������ΉpKϕO����������k�K֧�|��5y������>�x{��WYK��8q�����+w�iK.֬%��B�9J"S��ſ�U۸�ɔ��M�c4 AhP@����#c(Ӹl�4G���cU�2�� Ƒi����LC��sg[%�ey��L�8�آ���^&1�3��i�ـ
����_��M/L�y(+ /��"��)��U�^��:6������>6��?��ٝ��ܽ���K�X��!�ˀUY�6"�q١��:�/`^��W�v�Ϭz�c�kB���:"��z1��JP�}}��!(<���i�G���L�ݙ&��4��0n��1��M?��I��4���piW�X6�4hk���b��:���/x��C���Q�*�o��O<����B��t%�`���	��:� �B1�_���ק��{�mɿ�u���Ң�}����p�fNn`Њ��+:��gN�R�p��(%���.�d�܁c�D� e��CJ������G����n+Wiu�!K�la�u��n|1�̪r��K|v)E�f�.��A�\�Ǌ�S�������	˽w~�%���_�)���G���Bċ/��W�W������M9����U%<���N�:s�.�nF�Ξ���~G���^����c�Ʌ��t¶(~�Y��g��1��<~vg���?��h2ϪG�\�8s�;<1��I��k6�y�e�op@CSYy�[���C��}��۞����J7��S�3,�b���?f���W_91���q\K����#^z�?���s��~��d��h�f�	�*���S�`�P�r�����J�K�����V�Q>TL���`�޵�S\j3�P�+�`�H��%�g�)��+nۏ�s(�e߸;�kPv;1�a�ʖ�a�241�uyo�!:�G}���������8Z}\��?�4>9�o߾�p����#�%:X�b���iD<�&楤�����g�M�E!�iq�J��
O�j�O �H'c���.cM����ԕ��xJ��H�gG�9{������h~�)S��(�j�ٱ?Y�|���s��Av���"-�?����k�޹�y�:��w��f�/|�6�Y,�Xǅ����77Ǫ������
����`9��cé�2�l8vS�T|P. ¶s4|C�����B0�WAE�>�IC'z��pS��{0�?��h-��c�=g����M�S#Ri�K�y,3'��Ϝ�{H�3,�A�Z��7��C~�K�?���	m���H��z���v)�^�Q��n���QL�q���[��m"���uA�>�' +@Կ���Ð_������?pM�
��W�Et0|l�f5�͑�K�/�����c�?�ܳ/�L��I�S�=v�}���{0��}�Svyr,�/������WWjґL��<���X7���F��3x"_���tMX��ji�|��j>D�7<.���*��X>�iUex�9܎�75]V6o*l��P1�����&p�~aAR��������@�D���z9�����Lʅ;7�$�dN7��.�M��\���jN�Tbg�����?��#}C\[n@�T�'�2��͛7�-�wx=v�=���k�s�C��奕�_�9 �)a���!d<8�������\�����C!}:1�!�8��LU�@Vj��'Zr(�V%?	ߙ�R���t��S�p��5�I@Lr�[��dX�䳒�1�Ћ�5i�-�V,��D�dL2Pj(��]�@�!7�.l5�z�M  @ IDAT����������KCD�DoZ|���7�U��0�v�V&:��S�7o���q�؂!Y��3s�����Q G�윤g���� ��Avn9@���sl�$
�
g&R�ߴ; ��&*�W��R�S��.hJg׿���Ud^��N�Z$W���L0K��;�IQk�Ȧěd�vR��W��qx�����,
X�_M���4���p�	�o$�� ���zOK'��2.Ȃ ���8��8��u������s��p�&w�h��kx�Þ�Y��h��\�$�mu0A�^6~�A���W"��t������ʖ�:q����]��Ýt�����}��^��	&^�䊜�"�@����[K{�9ō�Oa�V��Ü����ɒڞx��d��$|��z��	�Adb�'��p���LI�|����j�MpM����
&�v\��, ��H�\��j�Oʂ��ǂcĦS��&�y����+�����4Ia��H��`S����	U=�["A��*��#�.�Lnf����w� IS"EG��x�.���-A��C�l�v3��a8B����{6Gૣ� 2��ɳ'�*���ZW06��<uO��r�	����dR�C���,%'ki���҃�U�A9?R:``iہ�L������9�5�ޠ����Xp<w�.����_��W���?�����1Ȟ8�>d�B2��x�#8U��a].����z��L�%�ɭ�(Q�,5G���Y7i&��#�J<e���=:(�)��ii��X��;��/�o�A:�·A-������N�\��&	�$eZ��vX��(��$vM2�$J�D�A!w]%�v�y��X"���`�0��r��H0�o���'ͫ���H�Ԫ�Ǫ.�)猀M)/��oU��^	+��`s���O/^�_�#�t�DW._��)S��#J44i�<`�^w�a(�3$5l���
���׆[K��bR>�.�oޗ�;W�ƛ��^�^ĸb%{��j`��]�� Y
�:�!%f�P��4K.���:���
�scC���*�S�i~�.�	��@��0�)J 1f;gSɚ����mP!UR>Ƴ���L����#��(r��)h���Bs����d��Ξ=��Dww!��2ĝ=����]�=5X��dGJ��O��Z��`��q���0�ps��*�|�a5��)�q�	�5�n�]�	�H�0D�B�/Ajv��� �)��\2���jp������A�<�7;�[p���l�&��{�|�˛��򡤯�a�USg��	P�z�9X��=�Iv�ɚ�(Z�-�H��PdY�����=�
$X���
�Ž�
�X� $���\�[6����7{R�*�C�K{F�!X5m�W�.����8���g���o�<��j,��ty��^4n�Y�KMd����(�J��* PT;��< L��B@��z�z�^�)@�d{diMO�Uf͚'�O���L�d��O)�������p>8�'=<�rb<�U�T	�)>1k-�vg L".�7��t���Ɍ�I$;U�>��;xVP>	B�/�`C�&V��ɘ��g	��'o�O�HO��Y 3�CA�R7�o�g��?��$IZ�?��T��a��S�?�Йo|�O�z뫜������!��U�����n.�B�y�N̻��" �*5� ݴKn^E�����=�żk[�5t��7m�o�Lb�}dS��hRD��" ~���Y���7���|�,A^7^��Vq�����Zb��.��MCW���OP�p`�6�;����v���r�e���� h��{��J��+A���M����wYhV;T=�*����|����叾��\��8g�A6J��zL�r������4@���������~�0-�j�;����n���\�̖��2��  �����G�4q
����L_qO��B� i}Gg����K]9	&;q��f�Һ�Zi©-�y��4-v�{�1MNHO�;�q�-���O}�n��&�� ��p`�[������|�|"�����`l?��������׿l�V�+!�x�Ǒ&��j�u� AT0���� s�extds��;:G��������_<�V�,�u �7ִIY����7�nCCG^�`�lh�G�V�n�,d ���Ѓk��3�Dq\G�+z(�q`��+i�.6xd��&�K�PS9�GNwO}\v�4����I�2�P��d#�ZsV��3ٳ%�^�J��� h�W*���edB?6���d6���kO>����EvG�9}�r�$���Dst�8�2c�W�pJ�P�1�!@fA�&��|����Tcy�~�@.f{I��5��@c*����V�� �AbhY��<��ȬIPΐPǺ+Wl���a�THJ�\nJw������z��󆢊�ܧG&	�S����G�GA��<2����O.W��JFnzF=��f���C�xu��x��~���  ҏ�M��Μ=��o����}���m���������8��ǥ��^�Uր �b�)�����;��a&���R��vaU���,I�!̇�`���w8��Jr���>,���/�@���|r��3hJ�,��-�̇ONGh�w@xP�Y�1K�W��Yp���^�CY�B�@��e�kY�O�����J��K9̙�	���p��c�=����/<�<��/���c����Y��e��2�=�G��H�LϜ:u�
��hY[Y��` n3͡ph�~�Ζ��X���Ď�ڰ��Uv�6^���nw��7i\��E�Tb�O��>n�KK�D��OϋH�Z�
��*�G�m$mZ+c����h���V�$ZR�5ٵ�G	U�Ki1� J��
���j֟V
�>Nq�?�3.t�u4�T��S1>�������Gy��GY���V��:����|�8.
?33���O}|����"3�|V�o����f$�M�vG������H��Κ4�8���#��P[��5l,0�%�"����)Q��9� gmY��D�I��]|J��[�<�� �_ۦ���&SǾ'W���,����t��� ���3`u���e��Ǜ�P���[�r�����R��@̫�l�f.���ƭ3�W�/�lh��0!I��ވ���嘛b�x��o~�/~�xNM��h%23�<q�d �~{�MRܛ�W�3�~������͑u����<���'d���e�ټ��HpiY��
�@p{ ��nCp���a"�U��߭Z�Sy�+�ɡY� }� ��$��Λ��dm�@I�?�3ϖ��V�d Rz��S�`����h���g��1*�G�w�>ZQ5�އ�N��+.o��;����Ϸ��$������lz�O�3�C*�`���H�s��~�iN��	����w���K��S�+s�4�s�P��� O�� ���n���zlf��H�'���'W		鞲���P���!�*9f�>'d����Z��թk��AB𡟜���j�ʏ�{)r��ef9Q�͆!#Z�rZ��Cd�XpL�r���NN�:y{�����y�{m�I^��e+��V���-����G��N6��]�u�J���*��4p2���b<Y��fr�Q�-xfL��<�!�LS�K��n���ѻ�}U�^U��� +s��y��Q/�]�=��T��S�[�l��9�˱��l���W�>���B13|�KK}#����m'�
��ر]W��&cb�v��<��e�����[7 ���Y�#v��0k
(�`�����jI&>:�n�O�g�֔bR����������\F�	��9On�0ϕ�����5Ca�V���B*�fg \��k�� A-��$�^ٞ���-7��	�����(�}=#A
��+�0��8ӗ�_�|�^�ɸՕDL�CI���.�.��	΅�b+���X�R	OP7!��+LQ:;sZ�흉�!c�#'����Q9[� 4}
�0	2M�n.W^��7,+mxon�t���:���o8�6�s�X6�s�w��n���,8&A}�q{�˯����q޺y�NS'Oqˢ>�Կ���wN�/�r� �)��q��&/�\#z(u�����Q]�ґ��9��;�	��l���2�1��g`�iX��d�6���zE��YŃ�Č��tn�����m<�n����y,8�j�̭LM������_|�y���׾4����/]��搕ť�����*�2���%e=⿜g�k����k�)e���X�a{[��՜hI��_W*NRw����%e��z.+��3�[D�M'vw�W�s.u�B�V)�,��|ڣ�C�)�������C�X��VA9�����E}������L�o��?�(���^��'?f�z�݃�|��^��َ���V~��(LX��X�ȋmGkl��wc=��캔�vPk
F�Og���rۈF�c��*Rn�<pz~Y(���.~Y,Р���Ydx�co�ęG��W �2[m�������GC�G'�_���EI2Ik1������z�?9[�(��J� �Xnc�.n2�!����or�����!�
Jy�	��>ד���C͑�͙�ӧO���T�c��O ��z�B�®X��)� !��3BB�����^��;���ŉ諐��c�l��諘�B9#!��>3�<����������^��舢��G+���:���r$���[��?E��5�Q`�Դ�ȺG�z�q�͆_�}��7n�do|�M�ĵ��R	� ��Q�<b=}����Qл1o��i�����1��NOO��r�B3��v����O=T���O�A��߼����X48v��*�9o��Փ@�`=�=L>eXZ�O���� Ќ���x�t�|B��wn��kPY�&���&��&!�	�8�f
�����?����׾��3OOL �.��<0+�'�O0w� l0�������Wp#2�إ�����׀��̈H����[?����ܻƬ�wj6Q7��
5��o��r�o�7�v���_�uOnyP
jN�{��>S�Uoə�ڄ�&Ы����Ӕn�O��ъ�	7���O�Xs�1_/���zN�H�8��6��P�q���i�Y^/3�\6"��+���䡝�g2�ɍ5N�aLcMb��I�. �"�V�W$��A�4�\7Y�3��m��(�G2jW.x�g���I �Ԓ���y��3<����T�W���Na�����B�y�ӷD�@��`ס�:�L[����Ј�}�;��o����(]�#:Y���Tn��.��/H%&���=�</^����d�nݲK�����u���]ǎcl3��Ѥ<�Wsމ� -��Ǿ��n��щ	�-��b�X�������>��h�3F�pLO�h0��p��_1@č����(ԗ�;�+|�'��r-EZ�W�$�G�GF���4S��������E�|zr���&��$�O�=�$s"�C�,�<`�k��R�ME䄣�yV7���R
E�Up{�?N�Q�l<�"c������L���:u��C6��Z��Uew�8���yT���܍�7Xa�r��̍�>[dW'��V��P�WWNLM��(�]�3Hm�Ɉ�N�9ۗɉ@}P�t�X�����B��=s��P�|�}��A���8���f~�o�YH3��l#z�gG�&�@ٵ�c���8SBv��ω�!��l�f��r�QGu>��M�B����O����������ǃ�1W�R�̹\�r���Э����9)�j�44JZ"��]|x����F�lM	/�& ���**nD��4�aNH�Fc�3�k��o�)Z���Ȥ��4kqʹ@Y�<H�T�fnR���i��!^���d��
��,I�Qe�����'�P$RvJ�	��M�4��hVC-/2��u�|{���e&�'��v��g�}��3/p�	�)�� �*s��=�jП����]��o{�ʕ���7~��,���ӧgW�u�X�����'�&�'5ʋ�ThUŊ�fځ%�4<��/�qP��y2"�Zb��y���� ���.\)fR�]�$��7�.wcɃ�Of�4�M��x�M@���W����NN��J5`� -Xx,*�P�1� d��R 87�QB�ikOhphJw�K��Ͱ9� FW�LNV�@�9.��Rr��.�)nՠ	���*-�'A$�
^
U�G�k8�;�x�G�Ѯ��2�1���P�X\���A�~��K�.�o.��h�{���µ�-N�Ff@���m�\�I�1��+}!'	8	MZ�/�����eL�d2�6�� S{`(������10�m:.h/B��Z��p ni�P%���6°�#h|�F�\�َ�h\��U����Vބp�=�(OO�۪�K�4�,��|�"Ý5�/�&tp��l'd����j=��&�؅��2�}y͹�_%
.�0X���φM���YUF�Q�G��t���An�j��2�"9GMV4�ȀW��d���T��̠D�R�gj�Q޶ͫY���	�";�(-��
O$��w��^
�xR��xJ_u��ǫ�rB]JiWpI*�pt|�V�;.��`�Y����ɩqzU,x�7b���m�b�#�9c���ӗ���yrCU0$]G����9 ���ȓ��'��GDʜ?Y"�.�*Lp�o�@i��&oh����9�M!Vǎ�ׯӉ��4���ʕO��;&m ��y�TM�঄��$��>'i>��t�E���㍈Ĕ������+v<A>� Ğ.��õ����A�G�.B���kk�
|���6��+|�Vg(n����:+Z�n[�vu6A.+���Nص}QN^K��m��m��R��o�E�A����W�[h�[��\EX���>^���"_�CC��wffN��/ I�!�o�թ}��(�0B۷���ef�>�-3�#��mi_Rz@����H����5�����Pļ(�|��܃��/z����m��5����6��J1�˰���D�����o�^Ώ�7��Q�Qґ�1U��a+-�8�����[��٦\��<q@��+j��*��/A�����I3����ƩQ�����t��C�,�H�wGUI���%����Y�$?��c.@������՛�2V�+J�d��*��K�-q�C�~�O���(:�qG5z��\�����%�����9<�|�9���v���c�_�o�`D��/hdQ���i`s�ے�՜@fU\��p�qm����[8�XqҜn����\F$�7*�<��:�n��E��8�pP(�%�a��'s���|��S�?2"����8����;�O�Β��1����M�&L���>���K�>Co��s��؈�-��h�X�r�5Z7SDu߅&�g7����~6��^|&l��rr��,�ryd3C"3Z��������	��.��"��t�+0h �c���`Ϊn�y͑���s��{~�����@f��ޏ��q!�T(����/������}�8FWR�HA,�,��FC*�N��|k�Ǝ�i]
���9ɮ��EY�U܊,0���6ֆo�dXp�����s�����C�v�<]�rbqֹ��:�lolWsO>�Rҗq�6�Q��.3'�薤.��sh��p[����?��Em��Ya<�+ZC}�/":!�%ԯ��GT��wO�^iq���M_���fN�檞$�ۯ�p\匫�O���+!L\����\_c����(�6���V�C�G�a�
�K_���Ìܘr����>d�r@#r��Me}%�kg}�N>�=	�<��4eJk�F��,�EP�-�"��'�H~�M�x�\����1pd|�n��v�4E�44�'P+�6O׮s{��S�9$9���ֆͫ�\W)�'nݔ���'�TP�i��ɱI*qlb�����Mf����ͷ�x�MM��>���1�8�kR��?��}�~��^󨪢��f�_���_X�k� �.�FpQ!ȭ���ǚ�g�͢em��E�a�Xu���J�Aԩ��Ƚ$A�#J�J�"�+azA��?�>�	��=�'�M�OZ6�o(f|����nj�ĥnа���������L[q ��?�h6�Z�����qL�� �[��V�5?a}K�p�u�,��ꏒ[��e����9�T7H�	ĀK�c�u�B�����ܜ���d��r�rՑgʿfK�&�����t#L�3p�gI���G�<�ڂOvdY#:%-3@j%Ȇv<�7��!ӎ�O�^�e�W������qj�����=�F/ćw;��_��hG6�ɾ��?���)��#U*Jv��[SS�y�%Ϻ���4-/����`��?^��f��)�vG�h�Rp�x�F�8�G���0�a�����9(�2M�zd����9��f5N�yF+��{���(g�?��/�������7����AHǱ�xxt�����g�'Ģ��!UoFѸ���s��ΐ���)�c@�:�3q��0j�;%ՀL*	`)��iD2�ɑ�~@ФD�6��^ ���U��P0����i��b�i��f2��e�b%�-�\�n��U2������%
ū��UG �_9&�)ꞔ��"��g�a������^x�y��B��>��Tw/\�ity;vk���w��ʆ�����׸����h��)��5�+��񿮀�Y'�3�:94�6k����{�S�I)�n�p�®J:�0���uG�� ح�v$�q3^�iG����H�ˊ���!]�����qd�X��3:0>9ͅH�<��h,1�}B�0���E�7^O�X5;-I��v}C#v
�0�J3@�x2ݚ���NC�S�*��$T;�����[��|����BI���t��ڛ�>�_�c�ʎ�����3�T���H�`�����q�REO�������ߴ�&ÎY:���v�iZ��iI@�¤�
�A�k���pA��_�]E��٩O`�ظa�wL3c�DS!�re����"v���&����{fv�nڕ�[�1��*"1j��i�Ǆ�Ae�휘>��|�ڧ\+Է��h�3}tzu�,�f+���6wt�PFa%Pm�i�S�c���ܶ��?Z�W_��Њ�Ъ�|D&5�r[�U+k��#�� 4����뢕f���Z���t
-�Rܚ�Z�9�"ח��LS𠫵�n����t��΁_j��>�	ARA��I��O�\�8��pܚ1����>��/�u��G�����������U�ff@3v�W��M��D�3�ͺ��fr�8�&���%��j%:�L��|�[:�C��r�6I�7����r9g��@�9�ٙ�Ǡ���P���`��d(ϰ�Bu��+�D�9�9�w�ao@���lj�9#^^�=SD���Gy�����k�4]~,��%���_3F�}�H�+�@|0�s����tv����*}���xБ����d����	9w�<�62*����öކ���|�{�� O�^���}�2��;d���F���z�Z��Z����'�������E��͖�\�X�l��XD�@q��e
��ɓ�3�n޼����Y%��weX1���i��`Ð�@�`��B�к�l'��SZ�Vs�!KC������fY2)��ɵ�U�n�ЋԳ��-��'�g��W���e]V�g�c�_�ٟ-#���iJ����EX>�?_f�zL�(��T��'�ن�w5Ν=˱�y��>��1�Y�`_:��o��#`�g~�S!hޘ+g�brr��}}�7�G]�*`��u����\&�y�鶺�{.���i�9�BH�jvu��(�O�\n�`��m�f� %�Mv��7�d_�WN �M�gh���:y�c����P��x�b�I�8���.[�؉�1������O8����}��L�v��=ʁ������LM�(�ׁ2V2 @����e͉#nXr�BL�Q�Ie ��^M�=�d�E�!��Oq�:��u�j&h��8c��~�.�B��לO�jѲ��9?94��y�i���
4[)i�2��$������p�'�|�ͯ�(66Fs:J�%�����ּ���i��ೳ3ss�p3��|�㶳�9���'�A�3XD:ԇ`w ��1��lZ_W��^QNv�+2�k�MR�z�r�0�.�߂c7��;8���;�m�:䧍F-h�PF�(�C8��׮]cc��������w���OpJ�U�1ḽ��	����:V�ݻ����~�&�t�X�Fc�����S���y�46�a?>Z�X�A稝l�WnD3@�x����M��4y���c>Υ|�¬C�`|Ή�Lۼ�����?�U����&Wjۜx��=�<����7����� (�5�bZ�B�ٞR��'xf�S��Z�pnnm���V��D������WTV�������UV:ku0$�'���c5��|p�5��H���+?����=ž͉���!����$3��}L8��`�����ի�o����O���8�A���5��TE\m����u[���V$}^���1�uO5׳�!��&�r�d���٫�ʈ2��%|�/��b����ҩ��K�XKP��ҁ�`��e�~�Ug�w֛�g�Zք=W�nmCyH[�i�f��VMΚ�����Y]%�-{E�N	�=Yn��r]��m�޽�/��6��7����H�x�8F����>���_��͛7/]��%�cc�'�O�+��O�:�����@��︢��7�iȚ.��I5q�hC��O�QN8�E���5�nB�@�� �g�P��)2 l��K��ޏʹ�,I��s�M������P��<��Q��X��\�X��c��f��s��ʏ��s ;�m�(��c�̏�X���S�{?.�	>�h�vtP)܍v��W�#�<(�� ���߼������`���FC�R�p(��c��9$�Y?[��}���	z��u��8��ޗD �c�\7��AF�^ّm�u8�<� �8(H��)��]�Y;��CKe�F�nZ�ƃd������R��$�0�<7��c�ӈ�P±wk(?ʧ5$�����@��|wG�h?T��x�s]������J�w��S��1"��[�׮}���˄����X�Á''p�����|o�|�ƥS߿cw�̌p^��f�F;	���J�	*��W<�N���^���	���#n���TIa��ACN<
��;HhuRw��RIA�z��6:Fo;+�#ʡ�YC%�$�(38���Ĉ������.g�y�ؽ�@�N�a�TN��&����>���"�6�gIӰ1�I9LNL��-�e��t?0�/M�޽w�"Q~ɝ�$q�Z�jăo)�8=f�&���j��Q4�5�o�F��d�'*[	g�V�u�������ID��b����@-��]>ǙӢ悞���C�E�Ld����Gy��Ϧ��)�TR�By���F���-}P	\���xfp�Bv+]�P�U��hÄx~�Y�?=����F*9(��r��rk'�]U�a��}sz�4�#;U[�,��R���|r�S.;x��s��C��Lԅ
AjTQ��p��pb�7���n�AT���{]����O:>�k�i�T`Ǉ�?ZAe��m�TF������	���b9O@��íG֚�5���ǁl9�!��p)y��q!&��
�̳|<V�[�͈��}Hj,�k���U�x���cz70�B���u���(�ч
ԃ>���}�n�F�v�N�|���Q���v31�2�'�&c���?04%��AV�?�s*����e٬9��_b~��Y6��Ǫ\e�s��4�u&�@Ã��A�L���d��B�l��MˋIf�1�����9�Q5�h���Y�$FҘ�����wM�<��!�l3�����z<��7S�����_B�m����sŃ��$��y�1�	�����¨������t������=���zq��f�}����������U��[�!��k�Ӑ�W'���)��$����$�K@�!�Cy"�"W�cui�c��{�9r�D��_���90pM�%[Vz(|�&���œW<������os��#,I�~�x|B�W#p~'�&�?�ơRC��`�ǃ#�?�K�&,���j��m�k�Ǯ�!\*��Ȣ`8��ޠ&����N|~�p�B��R�8��Z���ګ����(�H�t�m
_��d�S7��#�'�P�DX�tA��R>�<�S�����z����W͜�#��#���\�K��ެ�u�jI^�KU�6{h�� g&ھ���<���E8���1��C��v����{�Viiq{�6s�?�����Y{I]�����
�4'��^w��BT�k�IX��a�Q����Eś6�u@=j׷лP ԠK��m��<�&�A�<����;1�/b��zMݳh-��J�[=ͬ�Q���0_�J+J�cAO=��s_x.�5���(��%��;e��P�}�$���OFo7��M|w/C%�5���fVR��v����[wc�tL4MCu?�gDvS�`��)[!M����!({� �V[�[h}-n����Χ�oIs��5���釸�tzz�K����7	189BeL(��a��i�s��}x� @3�&5ܯ��ul��pQ� -��ʖ���6�I%]��*�LS�E1*p��	�_o$�V�	[�qȳvG�P�6��}��bB�(K�Ox�g�xbF{���,@d��48K)�}��g;*2 .�7� � wDS�Ca�D_�y����*�̬��sg�{����i[5�ޚ���?P{���կ�ᛷo��_ć���;\���N���`(J`&��Q2��ΔV�����·E��d�ɮ��Β?��vGf�;p��.�-A=���x����?�S��rgΩm��ɾ�'/�ޓ�O�b��,&ia[gal��[_��7�������4�+ 9�2Xoe~����L-q����N r��*���H1�ٛ�{`���d�4pUn�hhW��
H.U��.8"�U�^�L���m'�q^����8&�lY	�4�|�p@�\���n�t� ˙�@�n}��%��C�s0)�������"�[�M]��p=h3\��8A�l�̟��On����l�椺`�ª^tVDy�g�S��T�5�e,�h5�_�zꦜ�h��%�މ{��!��tK�U�kb���h����y._G�Jy�,����ϟ}�嗿�&��>���E^���������݃O>���f�p�ҕ��Q.�d�/�O����M��b�����l[Ӻ�"�R5ູM�we���מ�#���Kg���6��k�T�f;=d&�3wև�4�59�Iu��<Ϡ!�ps{X��#��{!����>�Ԧ(�BJ��3wW鶇u��I��z.kS]0�Ö�$��0'l����(��'�b�v||ʦ�������ˤ����<9��K/��{s�����iY�������Cq��t�w��5�\7b���;����v��зZ*��򷺀/ �!�C2^3[*5��;�{�	�t"�Y�����A��x�J�8��	��u�P�yU,�F��d��@�++ ��̍�~`8�%8yb�)�g�y�ôs�������A�n�j7��͓����Bw"1��.U-#X�y#�9Ɏ�L�m
�R(mڑ�e�cH�A�K���ꉸ�������4,ҩ�I���P2�-\:����\e�#����X�~��g^}�����[�n\��>	I��X�|=����E��a	2vꀀIƇ���d�#�IM#ș���j�������U�?ӻ�ќ󙱻{�vn���< ƨ�$9�aF��GFu���?��A���
�w���G�>r��-v����[YY�l��~V7��5?�-Fe�c�X���r@���Ǒ> ŀ��Qzy�M4Y�':P g�vg6w�ϸ���p�yv��h�<����~zaM�a]����a�ƫ��/`��A�G8�7���>�x����o���O��򫯼�����իW���_�-�b�~iiy��.��a���iF
�;��4�(�<?����g�GI����͙>�$�r����/v{�Vz��6�4�����	&�:��{����c2ǆ!J�)�O<�7W<��K�7�"h}ڔO��6c�a��5�([�1Z�����eA���6CK���<}p�d�^�Z@���ޝK���/�&�����#�1��3�E/�IHM�>���[[���sLC�ONlڤ=�?R���$�� jL�r��>�y�cKV�{<-Al����#�!S%����"R�`�鄰U�9��W����o�+t�`���w�����ǻF'NL�>G'�V7w��xߙٙ����܈�c��T$+�:�h;�u�M���/����9:���M�&�E���lI��Э�b� �J�����M��7i���eMs�vN�3��qw����M��䕋���R�Ϡ}�|�����1�鱮�+�����72$����g;�X�s�#���>Jflt�ĩ�G.<~��&'�t+�=�����������q8`lJK� �avw��bd~�^ce��Ƹj����!"ںȪ1������O�O2Y�Q������b�K�Y�c�n���\) m�cb����`�1fu��_���X����:���q$�$�2\�ӶAC	�mM�$���ND��y;l.�<4��o߾�_����+�s������p1�-ќ���@w��C�xa��N�M¨�y�6�/�W	�騨�j�@G*�2f��Q�mls;4sL�r>j�O�[�wN�_��N���9S���P��-�e��� �$�=v�4�E��	G~3��xRqJ�f��[bΔ���Ŵ[k�q��~ͭO���B����?|饗�b��rr*�r~8�c���kY�7iyy�����ŋX��2��		�g�=�<hF	�e�r	3>}}�S�~]e��k��d���A�xޗ �؈���Q�\'d*����� >5�V��I�N@,�uYw�-0��y}�mŇ)Il<��Z��b�W{X�s� zyy�l���;�>��Ͽ���A��ߡ^+����#���vn޺�����Nι�;�J1=9�>�u�8�d�	d;�[�d\Ճ�քS񓓺:���lx����#e�d�� 쌝���-U�=�O�|�'^ t�yq�Tz|=\���k�A��/�@�\�t��5�o��q�"��O�D��'���jc�c��|��>��r���>xeeY3q�He������x����|�	W�p�n����
�v��.*���&t-�x��7m�Di1���vd��\[h�:{�bTΤ�*�#t�R�§�[��C����h�z7�? u�h��B����o$D(FJ8=.��?@��&����X�)�Jr���yTe��CM9��D�A�6�����|�8F^��\f1�7���l��?=��5�k���K�o����C��>&{�1)��2C�s�yH��əH=�+u�Mv��`@-�����\�Xa��AO���l�`k9�������-�	Ɉ���H��r�>w��}���'�HA�k�㞨t:���F�@���<���݉���Qq�>�---0�E51�f�5��i�z�ai�:t ��/�Ȱ��r�'U�4����@�#&^s�8h��3�_�9�lEtZ �?��-��A��]I�h{?a���K��i�I�n�`���v��%	���P̴0�]|2}��̣1_K���p9ӷ𐮪��`騭��o�C�Q�l��~�:aSS��/��nn`cl-������:��iad e�Jw�LML� @��!�#�]��@9�4�4���O7nE\f�\���&�&���Op�W�T��l�՜����d0�J����I�����)	œ��5w�\;(��Z��I4v������!#�g�� p������i�4	m�ؔ4�e%�r�f�,'�m
D�ʎ�g���UB�ȳ�C�I�(|īƥ�����6��G��U��<�d8�Gո��H)<�D�ETߛ�:��A��B��T�}�rYk�@����!�2�QG&03l�����,�u�сQ�)8�u:Y��� 4��֯bc`p�"�����Q��2+��GW��sF����n7d�x5F�3�yb7W�H@���!��p縹v�GG\o*�k{e���SF
�:�h���xe���W�g!��T��ZI�  @ IDAT�y�P~��߾��\���1t/U��ɢ�4l;�&�0��K"V��qbt�_��0)s�����0�	*>WC�8�����Eӓ� ��0�ͣ�G�A��+EdM�qO۳G�t��T�g��In>KtO�����[�����p���5�Y��נQv�:w��+Y��i��=w�ڳfH�j՛�D?���cd�1Z�N��{^�:\�`!f��Y�N/��1P��-.Ӆ	n��a��^͗�`*F\���P�R�/C�?�o�0y�-"���н�2� �u5�Έ_2�Р��	�p�}
mx%��9�w6�6V�V��A
w_qsE������U�I�@���QR�OY".ECS����������w"��:>O#J�"`����jL'�̐ K�Z�	��[E�uƚy�A911A[}�Ϧq!$t�X���Ѝu ETBsw/~�JuG�G'?�g�������;�,9���u�g�=��`��\#vA�$� �i%��?���5I�I$�H����� 3�g]�]�xx��Ȭ���F���ٯ�ŋ�������7�BA+���R���+�i�ՅfVu�(�V��%J^�TW�x��X���u���[]^n�w��C����d�]�N�+=�E����>%�^�>�#��H�t�Z��ؼL�-����ݏ>���EFT��o4����[ñQXK��_������q�����~�h�ث�[c{��R�Z����
G�/z�^�G�.�RvF�0B��ɡ٤�\��{
M_&�G��y|jwb�	�8 2ņ�Sy[� �+�ѕ�9-������?���И�x"m�v��s)��ͅ���c���ݏF�)���>���eP�w�����e}yyU��Ɖ�:���`���[$+�E1^�Cz�`I�ݮ<s���]$��.l�o��`�/��02Y�q����� S5Q�>�ʳ���P��JT�F�6t8Z�~��q��=�&	Od7�=�=���_Xt���
��]~GZo�6����wQע�����r�\��(��ӎQF�d�š��N2�)c�lE�$���
ӓ� �Vp�:D�z��sM>�Z���"l�*/Cv�yk��yw�k��qrbii��C:B
/_�&|'7���xv~���0d��[Ʊl~���A��_j7*���ŭ��mzt��ؖ�X�,�1."x�zD�l*s-s��Α)K�!���-��'F��\u��~���֓i
Ȧ(IZo�	y�q�tF�p� u��݈��eȾ�5:sMjB����\��q4Gl
���6�<�^u�N~�L"ug�S��P<*P��q����s�lI�Q�	�[]�P�Id6���Z
�6�TD�F��ƧwF�<y�I�y㨒y+�o�FI� :F�76�B�@��(P��^(X~���N6R??�t�����u�����ĕg8�b��z�/{��v�G0�E ���z��y5�=�\IO!��Ќ��&$�i�4��|� 2P?6���-G��8귽�P���-���������}�I/!��u��
�}߃O*����?���t��z�L]�KW����`?��(> ��2p@#�hY�D9�Y��%
��5�B����/�+��a�o;i��?k��!� ��)�4qX��B��$n��I�}/��֯~k����Q�2 ���_!����7m>k-�}�<ڀ��@�X��#:�ޓ+��� ��ZD&4��`ݖ+Ző�	nb+���k��^���#$��o�ǿ�ohVZ�(�������Z�yYW!3l�!:l�.Xȧ�����>��/�^�M��-_x��"i��TKW-1�l&t@�^�L(ʊ����0���"��!��%�-*�����y%b���D%��ol2�^ l�OJ�g���)W8��wC��f����������q�����[M!�I�=3�dC�D3�����㣜�`� U���X�:=��O�,/��O��;��d~f�k���;���qy��Yp��_~���1�:d�BP2!�T;��Xĥ5[u���1&B��gwӾC�`��g)fĒ��|1�D�`MW!u1x�O*F��<F� b#~Zu���AB1�	�]p�A걶Y�'�!v�
����:��{����Lyt��I������Ç?����?��*�K�����BI�l�]�0-W�u�@*����ˋ��U��(>N�&Ĉ��w�K/VMf#��rQ�#�^�v~���s��[�4������������g����S�\��?�[\���Ŕ�������>������7�Z���l)8U����l�vC��УV"�_�Hۮ-S��볌x������.7d�2�v��$�o3@�i����+�
~�&f|�\���T$�"u�6� ��/���O>��?~�'���H�~.-�=f��Z�	X��u�n��gK����>���lEq��Ч�
c�[�R�5M�&(l�l1��d��J����S�}_^�d�#�I�-�K}���v0�&�i���J:v�Y���:-��X~NN8��;-h�x�Bќ��3P.��Qz5��|��M��%���'6�'�#>S�n L�?�jb�t���������������'�����G�X��0%g�T-ep��I+���j�� ��44������6^����o�؞��8��h���S�9G�!��j��vO�	�!p��o��&b��`4����0�,p=����� �8��y׈��]��& ���d�[}�P��F|� O�Į�){@�&��	1��q��ѥ����å�e�e�����{���2��ݽ�?�w��8����g?��?c"�ů�X��t��퐀y]YSu�T���/f�kEq�P1R���Us1z��ZP�,:�F�<��ۭ�w�K�30�g� 2a�BseA���`و����,V�uޛ���xD���(���.ީN������f��767g���}�h�y�/���*��\ϛ[�����6�-���ɟ��_��� ���,�j$*�ϥy�h��F��U�v�w�u�l����x�#R/�.�4���v�tj>J:J��nZGi�J��ؽ�S�:���I�R(��tC�q������ˆ��"K�9���d��u���s��[�c�UN�=L���~��:ΐ����蚢��%�GV�뭇�����Ǻ	��hYky8H��S		�c7S�M
|�V-�Ɗy�"B�!X��t����$D���rM�N�Z�Q�KPI۽A ̫��}��_�`"�pf�s���q�O��f��\���'�Nq䊝��i^q���9���a>�)tv����߱�Z�OFB6(wd���5�o	��Ҍ�{�hyi��X��lfvo{��p���q��p)���k�4g��$��ӟg�~Qc5aL}O-�ul&�3O�
�fw[V��ᙰ���� 8I��J\�u�ݖ�=����WE�p�9/��:?u��Z{H	��;3=M�o��̓0rL'�q���t��}q|��Ç+�O�|z�S��#�c���3��� tna���yY���k"g���=���	s��-,�}ն���S��i[W*`��	���h�i�ߤ�>���̌����I�g��r���[���|����`/*�4���t�]���:�W���̬7�P���'}	qj��hgg�������������d�C�����*G%Z������ͭ-�`J����98��SS�m-`�O����d��A��m!�#'7YW�Ħ�p�Gc�~n�h�2�i�@���@��ȸ-%A+T�&�b7 43���n(\��aI���o�ZʊR��l�7-�y��s-���8�!&vq�A����Ͽ?G���=z���
�g�?x�����8���l��{nd�����sӳ���a��q^}H{E��-b_�j����[pLٱvg�����2�ߣ4Id8=�[��lb|ʹ���3������w�F�7ɭ}rj&��sl-�++[�o�E��X;���I"�qE Ri��q��5�ѿ�0hS("��_�Zt�(O�|����Ԥ���>Q��k�����UԔ!�����͇@ӻ1pb����)���ǭo㽏��Q�x�՛�� �_�F�y����U�K�?>�������
Oulk�1;K���,	���~ռ*��+��Ժ�̔��,���8�uφ~߿)�J��Ģ��[�t�6�AS����4ΫD�M3!뢿��vw�I�'�t1��>)h��LU'7�	��8�Y*��#g�����n����ۙ����H} =dr��}���|�>���T�ԁ767�h2?3�I�rBf�[sX2�3�i'��B)ˊU��Nr��&5:s�������hH*4����0�[Pn��oH�a�����(\�/�d�_��3��ݡ��E�>���+&�0K�cc�G��pzl�d���G�7���ik�V������&v�Oo�qo(k�<�����f��j4������;< ���(�㩇�F�c�?��p��Pq"m��j����b�����!�Ws�=�<���F74�Pqz����� :�/;x!�fP�w�_�b}JO�dpxd���������+�jR�lݺ�wIwȸ���|�9�CՌ�,�=��=J[�;��	=>|Z�ɱ�C���͛#2��͜�)��@�J��2�i�f�G��z�?׷ʴ�N|�f�y���D���.��0��cV
�)���@ߣ� ԰܀C5�G/j_��2��]����l	�J:�0��q���@'��Zh�r�鶀��bK[��
�".>ǣw�Ι�ܙ9;�5?>=?:8����%g��Ll��4Հ6(�k��u���/d���*�\�S�����@��B��§ˠקR
�b�uI�F���j�ׇN����m��`&�1��D�e�#�l�0`	Y;��c�qd�`h�/% �Cj
7䎁Tc�d�[Mn�HE�PI�;�P6����8����FM�_o���n�"�YV�1�0�h�8�qsկb�(f�+>~���c1,8&���/<+F+Q��ˁ̼���B���q#��2~��2,-[g����ݽ=�������V/�8�3}rg�ԇ�Ƕ�Gfwώ�L�|$N{Q�NL�ơ�5�7�u8N32�-J#�y���|c���W���_�Y�[FZ	���h����¼K�`��c���o�v���E��mg(��<Xf�D�8sQ|���G��P�&e�I*�e�9�'��%���]�'�3�S>v�r�'L�z�Y�
� qs{ktzrl��q���{{juzn_�˼�t�H���X�РC裇�H���U���G�R�U���jN�5���Cʩ�b4���O��̈�#B�'�G�	^�G-����F�/�s����j�3A��".���FB����F�hH�-�yL�%C�7���5����I��.��� ����Ï��G's��NL�T�������E�.ad;���r��t�.d�⑫}E&�_�z�R��>�"gZ��m�`OVO�Nܻ�E��5��<uZ����oץe�5;Y�Ȝ�2g�G��y�5[�A�ϏA�ax��$�xm}�o���vA��0��@bЄW��S$�c����>8v��
�r�]Ǘ�Y�DN���΋�����$���9Uho��r
�J���'o���rr踜����W���-�<��&�1���ñ�ܡP�U�Z��q�!�3��V��r<���|8!շl�ký�6��rxO����Ɉ��n�x��*Wn��	�h��4g��H=���G5INSᠬC/ݿ�*|arza:K�5��9�����v��s&o��T8�q7��F9��f��=9����a�xu�޺��7�V��Z�ƍ�H����C"@"D�[�p�>���k�0�a�cl�-��5/k��9�C�����A�ÍׯU����ڋW�k��DG�����:�ue,�U�כ������G���~�������OY��4�4�B������9�aNm���N��ad���RV�ta�1���F�  �m2iR� ��T�`'F&m8	y}4�����`�/�����vƉȺ��S|o��<��3�
E�7�'�a��I|�&,u\�ԕ�� �!b�rr[&�����~�H����B�|*�=�B������8ф�B�f&`��}g�'�ci���\��u��_JW�q|C0�+�N[0��E�ȡ�9bJ⃧V%�i&�3�Z�5�R��A�����	)
c� ���u�ZQG��b̸@�2���<�n�/�yP�ctG�z�/����z1����&]�u	��&�N��8����.k�DH�ZK���F/Ư\i�ߴ��*��Ϟ>�Q�navG[�6;��9��y��(c�S��V�6 �y��iW;�Uq�с}&/��b�܄oZ��i�̲��a7oӁ6�j�b���P��=Q�>Z��������A�<����"Kq�,��cؓ�#�����[���������#{{{�>�Y�����[��IG�cK�E�Z	���X2*#��$�lG>I;Ig19�^�ڴ�~�u��u�HyC��N��i�v-�!�l�������Mܒ
��.�y:Q{<՛#���d�d�y/D�e��o�G�:iq�l����mml����>m	���+kkk�>!�u@BWԛz�u�q�6r��b1ozl|ogӝ_\8�ٵ��H �I��NhQ��Ãɉ���=X������_�@9�.Z�ܰv�Y����W�t�g,��cG�z���c��~j�i|��3ZS:�����H_�[�(@M\��S0�IW0\V��Ɠ�j�)� �a�y.�g�P(�������ۥ	�$����U��^wQ0��߽�7(.�J�z���Y�F��{�N�g�_ر��y�d���do���Oe�����dgk� �.Q��m�k�{�	\5��L��U���QOmjK����KL�b�ކ��&��5@�������O�T��d���õ�WZ�:5���� b@t�W��}.w�Ts�)����Ô��BW]o���qhF�,�v��>P��A�X5��1��(Q���x���ߣ��*\D8����h��+��	�d�2�����͔ӹ@�f=�d�f�:�L��!U{ì;pk����4��B��jER���C�q�3 ��r�c���R�EZLŁk����@8@ɵ?.]KJ�M֯��C�m�����7נ0	>0��&�s�P��ss#ӓ��N�X$�:��&r�мu8��h��[��9̢VVW[���bӌ�p�O���4>�F=:��S�Wu�<]�1GS��('���]��n|1�ů?�%� ��� $S'�$�0c��0Rnp(Hb������wCVn�`�6��z@}��w���S�Ð��"�bgw�����d+t�y\K�ݷ�-�����o�d���U7n��w����Uq��m��ŬB5a�)�&��	�B1a�WpB0�{�+Wۼ|���j@���	�-ܰ�����$c_O"U���c�̥F�'.	���|B��[���Y��q��Υ�2�ِ�OJW���9�nT�?W�~MU�᨜��J���/�_dLZܪ�,��M�{֞t9xO��^YX�U��G&F�ﭼ>���cb�>0�>�詅�a.��%���Ёk�~��DSi6���Bf{hl��;������^d`�`x���@�_>d�i���i��(��]$��]9rA�M�$^) 8�5�j�K���~l��K��
_ӯ�:���D�j�An�������o֪b�Hi���Aqo��6��m�.Ɛb���aEmccS]hf|���O|p�l��a�20d 릏��j�DvS��b4�����'���2�V�8�F+�o�-vI$���g8ka&�|������b�߮�\����Ҵ����֡�px�L]�O�n5��?�"���>��Ï��њ�QYa�U.�PU��y��D�DCF�e@���n�p@6T~�����;n���k(��:�|3��k1?+s�D��y$�t��ʓO����$����e��L����3���u�ڍ�K]NH[j�~�r��v}�!W�j�b�4)�����6��:�*�<hW���x�^�9�!r_l䱡�����$N,�9g����3YV��]E���eQ@lQJ\�K���rdt�ҷڇ}�.C���$؁ .���&t�9Щ���o�}=f_i#���&㦏&��ヮ5vrt:�;�����0ʃZ�hn�tG�uO@G_+r0�8GH���Ҥ3e��<1�x#4���JP
�ˠ���s��a?=�@at ��Dwq(`
'���Lt~e�
(�|��-w]�t�����6��	67a4���آ� s�������Dꃃ�ϟK1��q�׭ñ:Rzņ�2���6���V)�7����~�/	��/f^�̪,�m_*=�e��橑��+�xa2�y��'*�����Ĝ�>;>ff��h�ĳ�0u��H.��Q���3�&e�~{ѿ	�!���״=�j,��Q{H�]������8���Nf��[�:DH�m�7����o0��I�wtv���sSϲݤ����u��;S�΍^jMku�Z�`�O��[���j��������Z�ɓ'Z��3�[un���&� �8)1*HE��Y^�z�`��� d"x�횾Ds�Q�ڿv�s�@�i���;8�z+YI�ظ��4;oUfkw�8I1����:�{p�>�b+�1���#}�������nvU^��&�	�v=(Q�f�@+0\~-W[���/�'��_}I{�A�@��b��Yr�c�DvN,�RA���-{��1�͑�u���۫���G�3��}@�ݎQu*�)���Z\\x���7����E7l�}�ܜ���q�>��#VT�I5\�lL�N\����|�č%H��.�ƨ���;���ah�4����o��[0?��t�!?�wt�utp;^̑\�33�e��r�T�(Vs�U�Bīl�B��Υ+!�3Ȑ(�-+>�h�\!z؊���"��,ɌW��/R����(J�/��=����wB�q )tk.e���m��q$g���P4�����]���K���ش�g@���fV�y?��:}?���a����z���Я�؝�QǔR����%�g%A� s8��}�ɥ�XH�*�<hQ�7��@ԯ`�%��^�kX�ߴF˜ʶ�X��Dq���u�;�aÜ��Tv��$t��"�:�pЀu�2:a��gM��+�T䃲r����-M��N��9n/�xo�)���\g~nR5�	�`MR׋���.��?9k��J�)��c:�*�{��^�JG*d/|4�Tq�n��SӜ����M��\��*��x8q��@0��Q�Y3I���a��_�~��\�� @�������,�#n�_e��)'+�Iܴ��.n:�����tU�=�{/�q����	cƴj��-�vr������1�� Jß����}�J�g��P����7
�b��>�\�Az��c�Wj҈��J�^XvR���,_�"�;V��cN��V'G*`b0{&o>%�o����qxd9X��޷� ��~�c�����c�I���bJ1j	tvr��E��6�M�����Y�i�"� �&�����.����ܼ��S'G�Y��8�ޱ)� Hch��;�{{��c�X[�%^ӭb@�0�U���L�����'�0���~I*��(/�U)
��NF&�*6i���Dy_�.z�,�\'�YH�bR*�p_���&Yqb�QiqJS�D�lh%[WL�[����8�QH�K7c�0�1Ҋ̾��%�6�G�#�k㔑�{��Ӽ���#W=��h���v�a_fGQG��p1-x�$ID*&�r����C��鼋;�Ӿ�1n�8ԏ�ʡA�;���I?S�k~B��둃��s�0�Z�ytdg�h1�8�S�˰iē�A�����t��������ꌕ�ւm���8α������k7iY����5F���a�e/Fa�M�h�6^����sm8֋���q#��M68R."T t�/;P��\�����G����qOTZ�F����&�ePᰛ�}b�}��So~4#�����xĲ@jQ�&?Ƥj*�-� ������ ���ĭ��n�7RC3%@��2tF:M0��e��z��T�����.17�.T���`�%��n�?^��/�n��)���S���ή��6Զ�D����߻w�7!�T3N�'@s����7�xq\JN˶��5P��F��m}ggGMiU���f��4��S��Z���Z5!N�m���Ӑ�G�G�D9�H�'A��/ᶈ�az`J
.�����?K�!�x%��<�+3ܺ�#�P�3�V4hA�ͷ�h��&��-	��@VȨ�N�F���\�$�����Q�T��-{s�(�J�j��8�[3i��%�	_�9�-�q���Qe!���:��
p��f��9;��4��~���ވ�͝W�t�؛wL u�t�!ҕ(�BI<���+!/��:��u褃1{TK�]aZ��脵?|���9(V�r�blj�y��w���\�7���@�L�hߌ��V(d ��>Lf�Tt2�a�\)L�?����t�W"8(p����P�O���F��Y���B�J�j�#�j�c:��.�CG�84��{���q]uw�V���;�jb"&�h͓��5���pl��`gt�J�:b���ʌ���ub'B�?6j~�����Oh:P�c�@9�q�Q\R^dr:��P�����B�B�Qc���3���Xq��p�޾`W�y{��ʢ���������i#="t���<�!ƣ����=1����ufa�ܾ����c�ɩ�:������j��5���րpx�,i,��`�k�˒�;x���M~������b	�HGG|��k�.��:�<��W9�B�B{]DҤ�vÎ�b۸�{1~��E�Xlģ��22��3Er�!l#%��;�E�Ωb=�������������*�\	s�N��|3�
��ޑj ttd��rGj�Lc�9ɋ͞e]J���֘^���0�Y�C�b5+��T�:<bE�r$���@���w�>��e��".�$˗��m�O"�� �V�[���(�uܜ�a�]�I\�k�c ��pvP�K�j��i�S�0?쒭�лn�[͏���@����+8���1T�Zf|������Z�ӣ!&� b��{��h����R��Bp�T]�r�f�_ �]�+AO���rO�W�e����۽�u^��nJ�i�p�܎���WC��>VW>��	���̅�W(}NUd3��Z�02�x�p�X��h^nKP��z$�|��nɾ��B7&��\�+�q�)��5�a�A���	� ���(�T,�|�� �FxO���NRG����ܔ����fhr�`o?d����}�܄�����zK�a7~�q^,���`�92Yk��0��5�Un�GObYM��E-B�]C����2l.=6�H�1��V��I5�|D$4��%{+w�%J`�~ⱬ�w!�[c�Y@4K��"]��cLɅ�:Qku��*�`���[�HY��|������9��a��=\X�s���g��0���r�ql������!,m���g@Rs�����J�P;�%��W����|H�6�=��.z��az�4�Y��� �0�0 ����^�7l1)�J?�P�OM����w���-/X�1s��KV���y��BJ�C�+���/Y�d��x��{|���GgGomo���:z|.>jPL]�c��^�ї�VYqՋo�ǫ�7ʼ
�JFK
_��+W�y�Y=PU`ø;��sIZ
���cS1(	�GХ��4�jdrvft*�ǣ�㹻+�Z�R�եb}C�Z�ǚjyiɘl1/9�G���N<��9�@iZ��@��JQ�ַ6��Aፁ�|W��{T��0K��ٯ��u�C��+A�N�n���f��9�!�����G�n}E��؅��)�_7?����W���y��+:
=j�ի	�K�"H�~���JT���}��^֠A��ޮZ��x�+\Znb.h�X�K;D���x�Mw{bb=;��\���&j�6�'5�tN"l���r����搖� ��)(�������\~a�B� ��i��(�ΐ��n�@��6���嫫����ޞ=AZٗPh��<HϜ�-2ҍio	�0ʲ�g��1 ��'!Y�\�s�a��	'C��u�XZX���U�`����or�v��������{�����rr�@s9�D��͵sl�L��B��1�FK���k�H]3�l���?:��/W4��K�ë��ӸI+�k�6\=J� ��[B�%<rPj2��D�0d��D�jP���x+9Օ}�	�	e4�b���8���Z��C:D�56�z������6e�O����j��WWW4�ĩ0ԃ�=���L���*uE��8 �Tj��M|%����?�V����%b*�����/��|e�gЋ�ApΖ��x�(�Ej��`�����ɕ��0�Pqu��ȉ��,�m��D���:����R�]�z��ɩӄfF'�34?�#�/�^�ͷ�{�q����������%��{M�&ws��>�0M�w�lzڻ��YDmo~�F�X�`X��Q��E>ɸ9�ch����X�s/�K�eA��ۼ6>ҭ�58d�&:��cf�	�k&/�?�!���b�̓��cg�� I�Z��f[�cK{9j�4�l{{��t�p�(6~ǹ�>��A�97u�/j'-�%-T.����YY�f�z�3���X���+԰C���Б����Lj�u��6�[�s���������R¤<Í�s�4:!5���A�L�SBose���dx���DC�J�����������ގS�O���'�}�t�u�6��u��2�D�B�1?�����k�{ee���Ei�5�h���a�U�`����;�3�븃���- ݄�y7G���^������XUnrw�l�y��(_>�Lo'+�}�f��U)WM���ɴ��P0�����ٱ���E��z�fR�i�Un�w��P��&�S�6��n.�C�����|b\=���9�(rZ�L���$���<{��v>x@�129���|b�{lx#��p�q�XL,H�̅Iiv�/R�IF]t��j�͕�aH�J;��|����g9�ľ��KƘ͖���p�>�����A� =��v��c����PE��ǆ.c+Ʀ\[}��E�$�r��ܢtJ ����$u�W����Qo> �(#O��@�c�v�����q��qx�qy���s��|��:9G>&?~����',k''���T��b�!�8�a�7J�s""lQ�ƴIۆDf��"x֜�Q�V)ȵ ����@���!�oe#���n��#{�ܙn1��pH5IT����!�-b��-�(�� ���(���M���P�3ãm�8˃�����L�'|��ia~����r�<7�wǭ�ǋ+�*�h[��S��K�˫+u��X��Z�: ����"� �vEx�GO�����˺ťt�h�rq�2�B߈�דNm��j9�4+K]���S�����
�b&��]�t�Z~�Y�X�:��q���L?���>Vy.���z��[�㗯��H`]AY(�{}U�� ͆���7�a�"` y@L>����R���+�!���X����-������s�k]r�e�`�*���q�Ĵc�gM��|zLC�����5x������j;�)1���xz����XFd�9�K�o�5�F��]���1�o���'�Ӂ$vCth��L�
~=MV�z�3Y���2޸�b�QՆ�����X��+����	~�g����c�Ď!�Q_a��Xi�>l���;8qV1Fr��EQ��woɂ!%��R��7�kP\�fx �D9��sd@� �@FX-F��=��& %N�dJ�#��O`9����ȁ2ws��{I�Hꭣ*�0�e܎p\�I!��Rz��HHF��.���Ѣ!ȑou��`��z�'��8��MFO�N�f�}�t���z{����DH%Z܈d����l�d�B	+ZK���1�*:9o�H}�@;����%�11
���}uEg,� ��Cgs�17���γ��D�p�n�u�V��#b& ����"���a&a�M�C�>(Q��;���<"�R�X�S�2C6�$N�# ����$������
Ey�$��m�eltscciqqow'KY@QF5|��0:��=������a�9�"Q��3])3�h��߸EĪA��g�g��t�&X_�c�ɒ���S%4o��5h�h�S�&@�Cy��S��m`Ʊ��Q,�Bgl�9�s669F�DO�������~��` :���!��p�T�y��T���H��
�U��M�7oɏ}���M�eʆG��+Ā�'*�q1����`{�CU�t�rvw�8xmA�� ?�9[��@!<���4�\�?�894�;a�+Sg'V��ww���7��w���o��c�����:<ط��f��Nwv�
�<F��ll�	[{0�>Z(EF�&�تV��hI�,"�<�!2f0�2�X�u4!�$k82xn�]' aE�h�"Є����x�]���j@ܤ��؁�O�!ḫ,\������]�^�W�h��.��Q#-vX��]�k<��V��!��
��+��F���&N�N�6�X����g�M�H��~�Lf"���D�wt�᣽�����=c	wS=դ-Uy����{�N�:�=Q�?�`_��2�BXJ��#0�v�ki�
Y�����c7�o�g,�Am���3
5�:�D�Q�rӥh]k�u�7�+f�'p���6C��S��2rƩ�]O�������3��=�R�vxp��|bz�����څ�뭞rh�%���N�G;Օ���2�*�����Q�c�� �?l1�+��5d�"O���	b�yx�e�A"���d+�:ݐt�X�k��MMc�33S,�;{���&�<���OI�Wp�j~#��h@��a>H�hGK>`���n9���/�eT�cP����茲��y�S"M�K�8w�Zs5��t�Czb	�Di�� qpmI�'�MU�Nث��w��\���y�%�`��wv�_'�U��{������z_��.+�K��7�wU�	q�x�'��B��Z&Stsqb�1�`2 ���2A��3�FvvwL�1��AE���PiMM�5�	�{sI�ɀ<+��	���d	G�-e���xrP�+���&^��U�"ڿL4�ި(Q Kn�SLdsE:�6��"ᨤ�R����ؔD��*���ԝх�I�X�����������-\[=���|Ð��8�������Vm�<�){d�� )��{��k��_��8��[�v�a�E��3�#Z�/:ّ B��{Uݠ��q%�\���!�`�`-'9�4n5�⑱��C:�%�&�%� r�!eC���{� �P���S�ǢG��:=gp��'���9���daz���(��cE�_�_����ij�ƺ����iT00]'d��xa�ͅ�'t
�[i���d�Бq��%z����dO�}ysae���������������L���.ƽ^�+��7����{����G&(�o�����ա֭w�����'��<G�e�� qrxF�$˧0����8��2��q|�(t�e�� 2Cy�]Q�l� _�YBE���{n>քL���{X�,��nr�z�M���3in��2�C?5q:����af�fm;8q��5iO��{���1�hD�L(�hX�z�`2�<ъŶ�� 1@ο����ob�S�`\�ZK�h�r��N��G���P
�"��Lgb��Un�91��ai�/.t�z���+!�C�5�ƻ���,���	�Pɉæ�"�D�@Q7FS�6VW�Жn�ܼ�c�B��2��o�J��>i$JL���3�����8;���å����P�S��t��r����?�]�����|eI�;+�9	ƭ��9Jxl�&�Bٱ'��`(��dfrb�!)�Qv->1tٷ�:1�]X���P��k��A�0���ew�7?v��-DL�Z�:�a:d�2���c�V�2�j��d�Ɠ�-2��MD�u�7���ݝ���.d�I�5��s�n�X���Ȉz���>��r�!U1���0�|KX�����^���&�#l��>9�%_`tu�ƭ�a�8.Ѩ�.�˯l  @ IDAT3zksة��ׯ7�g�..kGnƦ�����ݻ<�f��v�F���M�G�㫌��(3�����W௄�Aa<%W�`MC�9�����@�P}��At�k��^ۜ�q���\�l2�A�H]�+j:�宁��,����6�e{{��62�6Pޑ�MEqP���~����UM�Ͻz���+���P�j�K���o�`��Pյ'��=��rń�7��L�Z�m��&�d�z^&V�Z��8�m�$�w��܂I%=9���1��f��3�sg���LQO�S~�PR#�p\�$�2}�f�f�I<K�n >�?�.|���������퉉8��!�(]}2�\������5X�Q�ջw��k�k�+�҈����|�^�Ӝ�v9���m�f8%W_
=Uy��b@���� (��A��ɀWꕁ���|�Ȑ!���Cؾ��9�������:1F�8� ����q���K\��k}mͬ�Qb�V��1����]�/|%l�������O �c�W�;(<�5נ0C����ܒ�>:�t��A̐s�&����VV������߿oS.o�R�v�[���ǏQ���>_���@�5m�s̺�5��6tw��n��ToJ�oÏ1
>㸭��F�����6�(z�K������`ɉ�+����/BY�A��j# �(������r���aƵ�ͫ��9tK�B>Bj,���_����1�B�C��5��cW���n��_��%������ި�Ȏ��00"����h���Զ]e�� 2�VBv|k�n��H������D�&����-���O.�v��Ǉ��Fb.�Cq4�~CxN")?��бv]¡m��;�ߊՖM=��r�뭯.ZQ
�Z��Ȳ��N�69E���Y�m)�c��Q��IU��II4�Z$`��v�3K"��wF���f�ά
��o���͜���/)_�~�fh0����j�B]ｋo]/�w�vzz������y�ȝ��9Cd2*̦*���8(�i~���)��rǖ���A@~��Yk��U��#U�eFg��1���5�	�޸���۷��X����>cG���	���f�gە
X�<�R�NM]�"� ��ZK~�F�@�|s�[�c�d����r�Z�~�{����e���
b�Š�����@8�A���+��1
t|B���.O��mb�Z]���������G�M[�o�4�7y�tu����=��QÉ�xCp�:���L�.�_u����������]�v���:lD�F���Ǌǻ�Q)�����.�V�Ɇ��?�����?fwh��t�˩	���=Q�
�l��|����C��N@,9EZXl3>��x'_ e}�"�
	�~�=�AD|	�1��o0�8Z^^Q|��7����툤*�ڸԵ�-̘u��o'A�gzAA��H40��y%n�N�E5K��u�&o���1�S�E�Ē�h�r�\P.#�8M�I�bɡ`����r��t�;O�=����	 ��&|�RH����J�C���H��Nq)5�d �th�j�r��Q��$�|p��鳉Q�8���L���7����ʖu���M{0�X^X4_�a�8ڱ��a��-��fJ0!���7F!J�U����ʆ��7
$K߫�\�--g�蝊=(�<��Ь
�P��8�8����X9�(�s<(z_�$*��f���`:�'�����`���=�,n-�UP�٣.4������2M	YmS�O�����yވ�_��C�q���o�2Ѐ���K�_���s�ͽ��_�-�v[�Sz�7:����z
@�xj.3��;�S�I��q����CO��|w���3>4%� :��kq�*�*[^Y�2���w��f�g�q�hd���q]���t���ݤ�/��-S���M��CBY;i%I4�8����ۣ�1��W4y�Ύ��x_�@��i��D����޳w�/��8��У+��.��6����2���hc\����p7��Ѳ�D�Z\���vM��:�&��J&�5���(24���l�[��O�Q�'��&��4[s�D6$�j��c#Q=<>�Rz�q�@��V%��FO���x�(",��|Ē�T�G��`�P��>�RE\M^_��̉�`������7>��;�W-�{�v���F3\�|�`��!@٩Df�I�F��T.��,�G�e!Z��^���J7���Q�y�I2�����rj�����xj�|�0TogK6̨����P���f|E􀡞���)BE����Ml���o�
���2k#�H��y�<�����.�A����������p�>�:��Duxo����k��%Sڊ�07o�R�֐Hj+M3�jjo�~s�5��xn]06���ϟS�u�Jb�D1���o�$����4�,����L�@���F�,����xjs���Yq�E=aPY
ݰ��j�T'w2z�x�N��j�rg������l�;�D�u�r�f�m��q+���X6u�r�2mM�JT�_�r(�z�,�M݆!�&�)"���	���W��V���̀�Q�r7|W����4�mç�u\���Z1o���W|}���Hl[*sb��gO3�~�m��rUw7��ɪ�͝M�4�
gw{'��r�S�_��"!"V����0N͜�J��M(M�A4�
�\�kSViBu�\�ʏ�T�K��e��C"G�d�`<�C��r���\�}�_�k��_D���=��p.hǁa����6�r��t���b?�3U�(��j�ͥ�H)2 ��飐���Ӿ��	���"�fG',�#���C_*��1~:ZV5���9��m�����
�Y�8��+����y�y�zTj0l��}Nu^�N�f���ۋ>�o|޴�[�a��C��̧���O�-�2�U���[�ѵ�K���Ѳ3 �h6F�J���;�c��s�	M��a	qxM٪�\��>��[��foM�#*������Ϟ?gӃ[8� ��%�ej`,��~�	߃W,J� ��~fHF_Ջ�]c��e��ˌc����\��=����@K�=������FS7��K���٢GD>��z�wT�����^���ګ2��1����}��}�q�j޻w�8�[
�f��\����BKᕢ|:�2A��2����3ƥ:WCD��.�N�^�)��R�S%���|Tf�M�%���\�۷q��u�3�2�/��D����NZ�6?�
!Y;�Z��O��h6DR��d������33����w��Rl������E�����r�B�#������DR��ڃ���r�0���Mv�e��P%��$�`� ����5�g8g�,[�o�JF����dAb�ŏ�6TKwB��0fA���N�����Uڌ\��2&��Or.�bl����Q��Hf&Yq#cbՊB^+yg5��LIC!2�������K�� 6,�����3��qzQ���lJ6�_D�˩�䣊�����ؤEm�X؁&I�T��I��]�J�v��Bpoo�L�B_�*��aS�`��DW�5��_1�̘�h#rH�ā�I]����Mh���VP"��KdqA@���3�����mwю}v�F��R�"�)E'H ����r���W���^��-�Ƕ���4~�x�ܰI`3[�r�����6}\16���G�N����l�G�4Lr9��<ZC0Q�c�����#d0�!.�-�L���d����D&�U]��oF[y�A%�{w�Mʆ�Xϓ,�\Ҋ�ʌ3�=�bņ�믿�ݡ���ސ���o3��|��ݖ��?N�GVTK���W/��?^�� S]���'jcK�ՂG��ڌ�0�K�7��I��ڕ!�L=�S����W�%QԌ��L)zH5�	M���y�<8^��:�WB�(5H��b&ޗHM�]ܷV>�}�ܧyU�/�R���R �a�����v��-ʩm�+��j�ȲB
�6�E�:"1s��Z��;1��e�L-��qO��x ����`�� A� 8��>�ߌ��8�6#T��� "6���Հ.
Vm�a����@��sC-b���B&�➗�A}\>ϞR����|��������ݖ�Unk'd=��=r$B�8����E\�q� �Y�{�p������ �s�q�����?"Wd�ߺ:pw<	��{V=YE��=m�
VS����y�����xy%����nX�pu`�L���z\�#�ӎI�GG�E��b -���vC�Q�5�P�@͘y�b^���Q�ѱG=~��3�
��v=����fv�v)���M�2��~2��;�a8ԭ'����Z�d85�Օ����P��͸��t��Ի)]�CZ�Y�V�|T�iV�VC�N-��L��ݲ���b��|F�u�n�;��t/��QU63'����͎�j���_1�zsil���c�ɾ"$�b��I�)�1��^h�I�-~��+��f�4� ���dW�iP��C-�9�URQ�;1�]i���K~��I�mmF��8��-L�t`zG�Y�%\v���R��}��Ի����]I�P|+�x��qee{s��������jm�P� �)�K�E�D�����3�M����xbԲ�7�br)*`����z���O��-wE���-�fN-�����.���Lh�e}%��]�q��4ԏ� ,�;"t�	#��]t�q� ���>W1j�ø���GР\�l����̫��qj��|�p��sdV��Q�E��yuUл���إ��WVV���N�D��lzKG��z=Rmq��A=�u��\��e�*�]��vX����0������2�z��@�@����:�A� n��m��1���>��o�f�Fg>(M�ϟHTGW�Gsq��S��
�Q��JVMķv���[��ވ�W`wuu��eL�R�����%�љ�]&����;��Tf8S0��L篦�㻥]y�M���nM���Aޯ����`�BWW���m����c���}eyACh�5�!�van5�K�F��W��3"g���b�|񌈦
��~y,�;�?��%�RtÌa�	ͯ�qی�gp��r7q/�;�[������	���j��>��$��"RS`CL,�+N��j��<d�ی�k��
�9&���8L#(t���hv-/��G�2x��C�@W�E�໱�(t[��d:��K�T�|����$�zjM0w>&w5|h��,!�X,���!3GA'7ޕM����=/n�Y����k�P�Y$�3�rhA �6W�*����M� �(��)L��?��):x��<DN�^&Rq}ٸ�:؎�n��8�9[�9���UK�6�8���b�e����֮���%f��n��B�Y��Q\`��b�V�P�$�t���R'Q�xgL������\!����WuÓ(ѣ�8��W%r��cW� Y�nf#̒�2խ��ތ�
�]oz��jg^U�i� ���?�P����x\6�����PM���lv���Şul�^�QN3�����3�=E2�w�\�v��\3_=�{�U\�:�o}�~r���0VWW�@�&|���\3�w'���&�~<�T�W�mԿ3�C�e|m��m�IN�@�/F�T�6�>i����)WP<;eB�	/]�΋����X�ߘ[k��R�s!��x\��/����z#_�3S�>OHD�x�����w��g���Y�G�dvjڙ�w���[ϣ��+��[��,R�A0%��j ��D�	��荀|��߹�� qYa�������5"�P�a�~߿��V��MLM�0؍��9�(sR��kxe��$�A�)vdR��t��N��^M	M�2��D�TWH�FeDҥ"Dv�&|-������Q�R�T<m4������T��|gznj�p�T��������G}���~o&>�*є5�&�ww����=����������T�C���������Dm�t�f�`@Ӽ�܁��l&GO�A7�:;ڹ�9Y*�Λ�T�:��ե��l��S��`L|=y��9.�����X��o�8�?��?�Β�6m5��d��rkq�ʣ63����>������Ks���Ս�V�UY�g�G��GW���	 b5�Z[u����L�f:�I��ѡ&��G�.�(��M�ZE/-Z��Zz� ��F����o�q��&GF�{����V�q����;K�sƺ0\q�������g?��g%�M��ێcY'���[XX�����85�V���]z��Y�)-4�X����{ފ����-�oB�G����̒8(W��0)W���?:�X�7];qQn��I�txUoSf	v������23��,?�����O��`�7����Y>�ZMqjy��?��?��/��0�Hz8f(�E�� C�o9dl"�6�J�ܑ�J�����X0G��ބ��`ř�W#T +:��L�V���<>��6����Lf027���M\H��=��+U��up��('��/��������z�Y�Vb�� F3�sRJT��5���Q]�&X��h��X�9j�f3�X@O���m��_]������g�O>���~������V�?����եI'��:2N����Q��㖹h��>��2p��s��䵚)`�=k9��C�&z�C3� �^ϫ�Q���|G���Ƀ+	��˓ �ٵ;c�i��c�OE�)h��a���;={t���~�?�яh*��g���	��ryv��v`]_��u���qmZ���?��������W�[��m���Ь9N��VD����X2kЩ5���	�3���L�
]�`N��nmD�KY\'�	�C6�'��X�^�$սa_Y��*����^���ʣo��6t@�N��C@C�3�hu����������?��̼�6��Ⱦ=d]a�0���kyu��>���������@����ݝ�S��p06���X&atX�*��w�m_�XHC<�oUoڇ�Yb;�ς�)`��=Alަ3�P�+%��-M�H!���zt�{j�N!����F�q��l<9�q[�h1���V���������|����rɀ[wڞں��������>}��W_}���}����8�,>������p�J�Z�n!��h��4j�݀�`� ʍP�ߐ���\�/:b���
�)��|ٗ�|���dd���D��e�K������ ��DG&:G�,�}!�vv�5/��d��n�?�TKGw#���!Iګgɝ,�/؞�������?�������r���M�w.C&����}gj�B���>*��W�W����W�Ћ/b����too��ɥ۾��%�u�tp���3ڣ}��F��֊�+0�Z	G�A��<���+�Ǽ���6�PL��)H�S.����S�q�8h��u4�V����ϣ�J7k�]	Q��/HOw8.B����q_�q����������?��g���~򓟬�{�zj:&1e+8�U�jw��n��~�u����ӟ�t}�տ�w�N=�����6y�h��������M�"������Nhvl;�)|���R�Ϊ�����-�$(G�V��Wv�Yx��5��b'�}ð]J��􁡄��6��I�Du���Z6$@E:����ah�bx�ti��>#��}���eG13��KD�Xa,id>��n��;���g�:���KC��O��lL���S5*������ȯ�ӳ�LI4C�*���l+h�����z4��J�J��;R�K�J��#W\��{x���I��Ѹ�����܋,����F1��tFlVV?����G�?y�D����9',�����N?i�9ǰM{s9�@������t6�_�������?����h�7�x����Z͢����a�l� �1�|]�Ч�':����fi�
$�ּC.DG���0�&C^����y|؆�:�96���X=%ex���zܯ�0|�.t���ÈX���Y�o��O�H�Z�0�6aR��Ey3bpP�X��lF��'��P����q�]I.��H��ɼ�ʾ��$���<�k������Ē������~j�.���43 ӃŅ8ʍ�I���I{�ץ*����s��I�t�������_�_ϟ=ǃ�yogKKqï�_ͣ��\ [JYe4S(>��A�vS�_d;m����Φ�bBH%���w�WN�.�����l���M�?L5�|���7t���Cʫ�bQ�R���1T�L�2w�B��f���[�k,q�a,���;W��ډ��� zoo�p��	A}�E� ����s]H���'�{���9�>|���#5�\��Rg�!2=��oߤ�<f�9��qܮ�޿�0P���x�j���g_~��/Q�����`fИGaǁ5m�����u�1/�s]X}u���ĄS51���A��ˬ3���{�V����F�����ិ�Ҩ��G��v9/5i�~|&�PU��S�j�/���!R�
���X\*�z����
�o6�����ߵ����w�}CH�E���ʎc���#J
HB�e͒E��w�+*Y��>6&���ңB݆ޱ�r7�Z��G���!.��ƐXM��w^��ۿ� L�5C0�YX���N֯^>o����&�]���3���9h|���B3k$,C^YYy���1'`���AZ{�Ӈd�����8fƓ��@YB�R���t�o�V��
�#�0���r��*5��Aߎq̒\�Μj0!����I�K�Rj��]4	&H(K��飇�S�
�b+����5�w�̆_ol�/N[???w����a��}�=|�#�=��Aoy���������^�)⿟�X���:���l*����uHraF���o�\�#�|���:@<{����W���ū����v�ono����` bo6l}��'?�ɟ4��o�������k_}�%}���G ��К�C����l��M_�*�Z�pH0�i�G'�]*���m?��D�L>
1D^��ձe�4���0��Ɔ���.@����}�dI-d��UJoI�o2,gR&iXo#-؃��yU�C}y���o}dȞD��n�Z}�����U��\.���>x�@�0��T�h�Q�4��~�P>�j�k(s�	���T�<��I3�h��"��D7��?���o���0��~��ۍ�ͭ�5@��XLt6_�B��w>�TC��G�0��)mK�ۿ��_�򗦕N������_����������_�w˹�0�Ƃ��(�<�쵊)��]���][��]YY��"2?5����`����YSI�q^6��Kn�riy�l@���� �6'y�5CD��*�������oVW����!#!g��on9�^W�v��Ï��Hn^Z��X�pl�x��I�G��'O��q�	�w�Y�j+�c�.����nA��!88�x�����}�[�υ2�~������>|�������Ȼ��469�{��ZW��?ǥ>|��z{c-�N<@���[ub�k��~��������͓��X��(Cȝb�����z����/3�)@o$c���`1$��|�����yy�K|gg;X��N�����f��V�,Ы�g+�w_�z�������˵�u#R�� ��x�����nnoa�^�<=:��~����X�+?H�C��������s����K���A,���p̊EE��G�Ϣ�
{PL�%�b�%}�����Kb��Ϟmq�/�����U���-օBzz&5�����G�^�I4iS�/~��F�c &��vF���t]hz+9��ed j��|�����1`$���_}��H�I�]�a��O�#?,�|Q�1!)����� TBD&Y�օ��g����qk���D�R䵵5�?8:����[��G�|�����ۧf�Ia~�-+Y�,D�bp��0J%�:=(�:�۾��T?����o�Tp���8e��x--�Z���/v��9=�)�j{cЀ� ��2.�K6�j���|�,���z_i��o����?����W����~=51��o�����P�7�<;=�#@`k*��\fZ.�z���4	>�b�3����sk��������x�l�`e��	��;�v9�N���;=>��=t��A�L�}7�	��$���]���ugtllny�]���O��H��7����㏾��[ye �dޑ+,�󋚗|�� $�;��Uk�)2�c`w�.�Txu�i]^�L��9=����8O����	����~����ӧ��?��?�����_��7�-�B��2��ʼY���.$}��)C�����c�@Cb���&�եe\�'��y��#9!�RKB�M(<|��H���/#��&v:��e���}�{k�ք�<yCD�����r�(_�Tk�k����j��D��}^M���D�OZ��qH]�I҆�������iʊ�r��b%����8\���;!x��#1S��Xڃ��=~��<P�� 
"R�OC{��������R�3�a����u���j"������*�c8⫵ ��C�ÕS>tι�0�;�?8z��dwg�^l�޲���ܜ"��Z_��1;?O2�P�1,� ����g�tO`*{�e]������]���vO��;]�����w��7��`G������*-��P�F��8�j���Ez繅E�?���`fO���u�������@�/掎�o�eQb�[�@ˍ>�"uX1��[>$uJ��8�+�󳗯�Sꭿ�0�%Y�x��!��K���|���+�t�`�hV`� n
DZE2�.vwe�%�a�l��ʊB�Zn�8�&.�����j�o�87~�z��x$�%㬜�Cwس�O�YzȑZ�`7���9;:?s��9I�%�6ßA3�cӣ��U]X�?��o��o��կ�z�<�0����X��/L�Y5�K�/��a
{w��P�b�N�LT�ʦ��-^9lN���8%���=e~y�>��	��C3T~����4#�++̉'&���ķWB��/3����]]^�����͹�i��+���a���c�S��39[��g���>�e��pw/d]8*��k�?u)���UG�N���S��A:���'�vVzc���O�n	s�y��8(��T.�qCg@�(���|f눤:��W0"���~.���Z �yL��M<+�#�Op�&@:HH�G׆Z�t�}�ᇔb��r>j�*?|��=!�������}i�4M+eqai1�壣�K ˌ�_-�H(k e���-ѽO�c�7W��j�2�;���$�E��{W�^;�[N0�O�O'���n�|��|	@F�v�UN|O�����c����)cy�0}��鯾�����vFs�1�2U*��D��Y���O��m�� ��	C�Lc�1#i�v~����@+F�3KqqJ���K4�>|�O��Og��V���E�o��89<9;<�8�[Z�!�'B�%�CK�XLV�����#AFGxb���>OU;'��33�9�V�56RQE�gt�EY�����@Ź����5����T������IZ��� � ����_�WH��a�{�|�`�&��cM�Ꮕ4I�׿��`f�hr �\5�t'WƬ?N�$����? "
)%iJ��99a�1ny� ci��'���v���!9dz.�o��{XȈ�B����O��	���B�}:c����T��(�οZ_[���ἡ����	��Iy������,f�^����Se�������*���Q┋V�h0-h}�;��o�{��� �a�]�� R���`�[�@��\�焏��I�ĳQ�Ѣ�vL���9|��O>Y�{W�'��R*U_>��
5��,��	��%�<1H����c�3֮`�����Ё���+�E�L���������/���W ��(��\�d�`�\G�g�dka�0�2���U����W�I��oC�N����rD-��v�.;3�����+:<����W��BKG%�c��~�>S~|7QB0?��'Ί���\��m��/�p&
��o`䱄X@� J(�Uf�'�/�I���7B�~% *ho���0T�_�u�"X���1Z���^?x(��!���"F[��3��g�r<ۚ|�U��M�U��1�v���u�^�ؼ��	�F�Ņ%e�h�xT�9���~��5�q���u H3{�5�b���_�	�`�6�,��	�Vk�Wx-�5�PB�FH 팣���\�H��(�>��L�����o���/,A+9���J䤟�}�viv��������	�'�G癚
�<3�rk�̌hwm��`��ʴ0�!��V��C���+��Nd����R��o���ǭ�Muk����Pa�X��u��N���9(��ҟ�xP�1Џ���4 &7xs(X]nm۩WY����(*BF�+��;��0��$���U4G�aCM��cdg 9�|��ǔ}��:�5�/�+������ǺbHE(��ؠ�����
Fg��97�]5 V�n�&�PF'�x.�n�s��]f�b��S�k����}S��Cg��!b��T1c7�;��[�vTsll/��Nj<�@�/~��@�P���f�� P�C1WVnA!�dqt�O?����;���ڢpAD�~ٰ�3�B��� ��Es�(I$��HJ������U�"�a������O��vsX�ُR��S�csӳ��ŕ�����!��6������}�IS���KF�^l��r�TQ�Ŝ�a����z�-�Mc�4Ц�^)��b��_�f��{w���q�� O�D]�,9r9�?p�x*���c[v*����$H���wHRd;�K,�J�����;=�o���↶�l�F���T�8;��7)�O	BvTݺq�3��\��ʇ�O�w��g?ݽ{���1�oUv�v��he��z�pBd0 ���U�l6"u��{�:�*���e!��t.7�&�0��nc�x0�!c��`O��&lP�]��2:��rUN�k�QZ&��Kdp�\6 tq�UF��4l���;� ���~����注���Zr��-�+{�pq��K�ѶE����C	�{�� \�.�zNϞ?�ٓ�d,���ee4q�����_��m,����lF9y�PA�&����t���b8KUʤvHnzyJRJ��R`�g�K=H�oְD)�@Y�T�sDA�;;[85�`�y��_z!�E8�h�T@��b���V?@���2���~��=ە���5�c6.%&�����->?-�l,��]]i���ï����vQA
�����P�%F`y,���ַ�+"��H�~�p�Zi��)���8�Ǐ�ov��Ȓ�Uբ������Q��`���L���
z�O���_G�6 ������p��E��-yl �и0zyfM7��N};uR��cv@O݁zU�-����K�]����B�p�<�'�D��X$ٷw�ד���GM3���O;������^z�۶��	�%��2ٗ�,%&6�bl'H��Nt��Hb�,�x7�)+����EcPN�X��������R'`4Yu�7�����C%e ")�r�F��KҖ`N��1K�����O�l�d������4�{k++��^c��k(y�r�>7���{���;��߭E�\��?n4��5Z��ظ�Nz��'kM�B������df�sO��:�M�]m��w�������h}���>��?�!p�)^����%���W�$�D�S��I9j]��;�#�4�=��"$�	��w��ץ:Lӎ���B��W��^U|2�035%2!b� ��5m�P����?���Hc.766N�q0{-|ˉ�5�G拠M������=�:w9�ֈy~>�7�Χ��������fee%�;��_���T�퓞������Mn�7��b�x�^�I���@|yh�e��>�/�3@�2����ki�/V���kg�`/��\'ς2��8$r��b�M^��66DQF䤖i�A\���R���g�5:aڶW֠6[��$,1&���5�]�5D?床�\�OM���K��;��c[����n�(��<�fC��M��B�00P�B��|�f
G.`1*YS��Er;����}	;,g����J���$ �^�[$����k��l1���������1f�T&A�cw�A�9�+>�}��Wߠ��W֕b	�8�儡�I��yW�y����|�_���I$��/20NN�)"跷w��X�X�����J%Mm�N�^$��~X��a|��c#2q��Ґ��c�\���H��Q<�i���P>��"��H��f&g�ƻ8�Iw{�h�4�Н��g�I�i?�j�[c�j.����[�Ğ�����G��y�	���q*`�0�b(��D��n�Ɣ�!.�M�4�̓T�����os3Sk�K�ÓC �qB�d����$�"��1����O!�D�������*�
����#C�@a��D�	�sN���u��f�x�K7��̐X5��}������761�K���GE���nF(2����&3 ��na�ǧcCÖ�%bU¢*O��)i 
�:R�gtdL�I�)&�8��q�����ж��l�_��\��i�D���=3s�>~8c�OVH��밁g�	�g1�ҝ���� .��F:��$��E����ϗ��$��4e��u�M��s�����O�������$$Q��	J�S66֨#��܈���$�dK���n�ƒ`	��'��Qț4J����+��tlVv�F��#��.���X��_�P�er�{�Q77��+�@�4�����i�cP��U�zt������<�^�Ne�<a�gk#e��i�E*P1S�
��Y��o�ŝ��w������0��5�K��'���{䛜j�w����NzRK$Y1����q4�gϞU*Ux�pzz<7?�]bC'�Ѝ����ܢ�PN�;;vWP��`�RF,P�i�hou� 7�a���l�on�|X��Q��0(��\}�[B*�c`ff�յ��&�ǰ���\����Zc�/����;�::8n���P��v�iq���351�:��X�5P&�E;�s|�$���1�����Q^��\{���CfkV\��2� I�$��5�nm�N�aiiI�-9qy{[����e"���S��/t�b�1���F�'*�f�UWA���>S�m��������bO�
`�;��JC7�0��t	�S�-��i��q{ŏ�X7����㗷�Ð^�Y�F�{zz,.;& C�&���*u���������nno�/��olmƜ����)������(O����"e��ó�����9�����U�O1
�D��a�6~v���ɀ���f$fk�ͯ�IJ(=Co�3�-΢���W�֌Y�^|������̰���c2A�U�!܎(�4j5�oߺ3=6�*q��Դq��0��*ٖ��+#�/���mup��^{��Ȥz]~������2����g15)��EwNU���74��m�08Y��
�����9�	
��b�r�k��'L�����l��x���8�²5�^�����0��$.��j0�z w�� J��Y�k�s3�^y�:�->�C~�������
��WP3��t�Ν��ݻ9-׿oc�0*�|w���m����ѷn�7w��:$"F���Xb���D�꾁�u�'�O��N��,��_���f\�~����4�o��H�(�zD�L1��'������{Y���7�F�X#-K��4&����Fx9˷�ލ�٩iS�>&,��H�)�7Ч&s��OY9���B�	^�q&~zb|rƜs��#�<��65<Z(���͞�.����?��?���۷�ܷ�����nV<~�1 ��I>�ȕ�S���/�e����������-�k���Z[?��c���ޏ�dT	�A��h�i����1�@�<Z�)��K�h���E��<�٩(�7��|�*N`�B�zw"�Z�k$��r�g���'��]�
	�W�T�}�������!�~��M%-� +\\Oە`��^_މ_�_ɋ�8�5�c�Hq;�3��ř��Q ^O��;��|�����ʒ�X� ;cm�@��ǡ�f����rβ#���1Z��{��F��>�C�M�^�@�$��MY�b���s����Q|M 2#�������F��3�i�q�!ܹ{���rX>}���LNMR�����Ցǯ=��cx�"u`��  )IDAT֘t���(�ӌI<�o�}��j���K��fr����
�aG���T4�m�eʯ_���v�r�2@������;�&DmO���pM��J\5��~��&�rP��6>�0��sΥ�F���܍J���4:bvv��v��X^��������T0�Eߑb���g�-̨����Uf<q�)���(���T�*�hx�d/{/�y�;0�xI�`�%�Y&	dmh���6��
{�>���f ������ӧLFWw]r��B��I�r��D<>)��	�H4�ۭ[�t������V�Z�{��F�T������7<�K��.����ݽ�X�˒�N J����Q;ums�Y�1F��%�1�gD����/cdd��]��|r<���3��O�5��-�DE���(���)n�o>�t���f���@#(�i��n�(�c|��*�*�׶ܻwς�C�:G5�w]����-���<~~C����~P����K������b]�V�ג������E���z��t��H�g)Omc#�� �Q��#׉R�b��t �Ӊ�I�������h楥%2�puQФ��1Q�;ފ�޵,�_�=7!>[ �N�g��d��7hk�J7;��'ow;�ݮ���#CT�TL�#C��ZM��E��V,��,��E�Bz��i�;����K	&#��\�/,�m�	��<�ɘ�����X���\ƲJ�O�<����o!��G"��V�=k��|��۞�V���+D����o�o���O"~Z��.W���d�P�6�3K�Dq����)�h� �P����wP;<�C��*<�L\�������9���7�f_����M��<�ٗH�H�k���;ۺq���P���^�����Wd4�CW���X1`�j��ha7I�lS4��H��γ�k.�-ЛS�����P_"�g�Ia� ��i�t�:i8�l4e�+J���tw�ūo�z?>�O	C�?;���=?���l:��e&�Nio�g��j�7�ёǿ���,5�A�/��?���m��w.;��{���6G;%\n�����S���u����x����    IEND�B`�PK   ��W��s�2�  |�  /   images/fb2015a8-ad74-4a61-8d66-2e77d7201afb.jpg�w<���>��V)E��Qj���N��:���*jDR[�ԮZmժ��[��gQD�P���g|��?�?������z��}]����:�����I�u~	 �� d  �Y�:n �i�����`�w ���߶���� ����Hg �ǜ��o������3  �O[�J׮)'���MG� ��?畕�>���?��όtC��w��og�;������?��������?���� � t����@OO���p
F&���ӿq�`�7��,��_MO�xz��a:����?��^��
�:h�b��s�1p��:龞j|��X�?F��yj�Y�s���t�L������F.&���7�\0�g��������6��x	��oBX�]���$yEJ������������w��=|�����S��/�^9�x���������GDF��NLJNIM����k��¢��U�5�u���]ݘ�=�#�c��S�������յ����߃�#��	�������zFFF��CG���N.F���g�o�3�{]�|��f�6q�x��o��]�P�J��ҿ=��P��/��ס���6`c�;]0. @]�����Q�3�f�t�S��N�O+�鿢� �Lt-3YȘp�K{�(��
7T�~{Ra��W;�Q����h��lt�0��r{�v�8�x��ېF�����w�wam"�;Į^��ɬF�Ã�:�Y/��s���SQE�Q���ZZa�J�m0��/O~� $�I�W�c0�r��S�S�jT��M'�[׸��kp�5�r'ʸ��w8}�q��'�hw*Ã�Ľi ��I4��83�%�1���.�|�[��g�wx���}���(?J�R^�E�B�'�(��W���M��t'��ľc���\_#t}/�+�Y�v�I�K�^�@B�:�p&>^4����9�N&nhCG�h���A@��%"2�$�(;��i�XX��"d�Œ-Q��o�l�r)��Y�h4���tv^�c,Ef��$�#�X�D����U06v��2j�?s���՗D���$�%�������8���A$�c%�J��7��hhRȨ����y>A$?����a���U��@�}N�o���v���d�!:��c��g�zX�fz��U��^s����jj���X�f�����b�9��z���H��<fN<��<�����%Yޘ�y�q�>�B�����%�ѠT(ȗP�<��Z4q=L��[FƩ�5�n<4�g������φ���S����^��1�"���wt�?�ň�,g��A���Zj�W/�LYJ  �$�e-/�c��뎮�76��8�\��n��N��gQ�[�-��y�iu�g�����Aj,*S���!Q�T�F��	��vo���:��q�)�ky������
��݇�7�_p�$�gܷ˾�)�y|�z�q��u�!U��UQ%��1$�R�"�.[)��\��&B�W��b	i>�ܙ�o�(u��rOdn�٧��߳w�G��]%3�� ڌbP��/C�b�C]����Y�����N$н���[�
FX�`TE���~Iĭ�Ǉ�f\�ߞD.xl~�`:*[c\�s�غ�6Қt�_x��]�ph�O�.޶���۝{;�Y�C�H�Y��9�K�fصNXj��qі���I��}Co���䑛\ϼm1�4�{ X�1�'�u+rC�7FTM���m��ϬX�5֧�ɋ�d� ~���+�C҉18��/C��+=q~�<o���ϔ�
�w�fi����Ż$WQ9�(���7=�[�i�$�cQ���slD��i�A��!��4b5�R���6j1�8��̊�i\Ņ	�ɯ��C*Qdم���h��X���/C�s����~#A?��*�PNT�@�����rD���&K��C�;��㾭׬�T}s��P�]�]��:�t���Cr�GJ����n�q?l�19����Kiv�W1F=ɚG����s�e)*؆|s}<�k^2sT���:��@�t����Z��!�aJ�v�%1��A�TWBQ�C.i�/<m �	�g#r_�	RG]�|���U��t���%/�uJ��8�Փ�R��}'���w|�������\:�ߔ_���������]��N󦐮<�;f��]kxd�V[1��m�['P_�Z��H��#%�xi�;y�E�Z/�aZ͕pK�9+�0��EM�m��v�X�0��VP���O8[��Q��V�
����F��g'��4 b���o�a�ߡ���K�x��Y���1�cã�WQ���Kd&B�0�ӌzq����[~�`�nvN����%n��Lq�C�C�S���/%���q=�z���Z�i���� fE~s��
^&����zw�`8�`�.}�������;Yd��W!q�!U�nrLF��r�L�d+2�R ��7vz�����s��W[�v^�����x0��?�����/�}�7P�]趭:D+ȅ:�m��^Ƿ�%�ձ�ݘc� �&,� m�#��1���BJS7��4;����B�[�9<}%�r�K�H�7��KQ�*-��Cc 	��S�U�1p>�� aψl���l�:�=LK��EbjR���R��MS���ˍ�]��A���Z�A��Gn��tdP��^��@b����ě�=�ЙxN#bSek,H��{�
��7�����K���$�1e5���Q�&�f��:-&j+��Cw�j����z0o�pB~��J��\A���U���R�x��q�Pyz�N�r���Le��2��U�)�{�|/E���P�OGT6wq�I$n���cgh�@ם�ɶJ}j�|\�v榰_ș.!�Z�h�)���f�t��Ker��+̶$sꨝH�id������Tk'����o"U>?��H)����T�[o���MT�p�i��L�&��'�1���i������0���RG/$��,���#8��Gy�s��W��խ��Y�녑g�|%�[ݙ��q��'������uCtN+;�d������Ӽ7����9	�}ش�CY���5֔��|�>]�$�}J0�Ńz	�U\�.-s�P��xR���1sRC�d����c��6u	!��g�My����/�kA�t�L�������ήW� ��u&d��M�ޔIw,쑵�F3LW�C�B����ݸ�A;۷�8�:,��EE=�/��Ň�a�\�F�'��fr��m~���wb0~q���I,-^��f,Y];�`�{�ȏL~���<q8�W��?\�y�j�/�n1�!�j�����O�~W�Mfd�`��н�f �C,�f�Uz=���݁O�C����tm/?6��>7B������g�c�J�N-8��u�a�2��ws�u��Wb�ʊ�H墎!�����A���5�y���R�Ȉ�lK�.JUۜ�?� �U�+���#�RU��cWy��܏�HZ�*�KN��ѯ��j�ڄ�@Q��|Z��`t���~�k��c͑2+�À�-���7_ͷ�{a��|��,um��ړ?���$���T4"�µ)�-��yb���k�v|���4����#rW�n��9S��O��B���G9�{a]�o)�ֱ����6E╘P�3�����+lc�[��Vw[u_<��+�ҵ���o�V��!xG;y���c1���S�,��޵��-�	����N�+2V�$�e@"�~g�-|uL�9���6�/����&|K�b�yk��>�1���;دS� gy�E�u�s���d��i�?X��ĀnF��Լ� ��
�/�;�����~�e���b"W#V��;��I�O�S�gp�{�HĪ�UjH�G��n:Zo-Bb�R�ٗ*�oH�����1���ϙ,����� �f[ŋSU�牛O[F}���|Y�ԽQ���%.qL����j"BJ����/F>S/�(�й+ ���VB,T<�Hu�2b�BH7�j0�\��DR�D��=Y+B~��ņ2&����^9��p�0\\�ſws�1H��&����\X}P���{���M�%W4Q����RVX��ǂ��(ǃm4�jѣG^9>q����B� �Y4��:� B��S���r���k�v��'?B�]״-�M,8١.��{����l�ĕۣ~���OW�"چl�EK��c/z|z.#����W�>�{�b���ؿf��PNӯ� ���B�Ƣ�{���b��],�� U-�׵P��5���d<��2��Y�ݏ�Hu�?���V�>߇S�����n����~�h�3'
���>�u~#&JR�bw��5�8PP�E����"u�����P�X ����6Hz1}�C�A���n��j���Л�8/���sT��oֵK?�A�/2(v�NvU�S>�8���:����s1r�7���������eO�q��I������>�h�Gx�BV���-���O+�q��]']�G�	7m�Il� H�S��7��ܬ��5v�yS6z+!�hCdob=��rѣs��8y?=�a��n_�=x�;$]*�/xM��Geo�dU�˞�E�ٺ��ҸZƺ���s����g�'��N���f�>HZ`7��#����wܾ�-F�5Lnu��v�)��G� Y��~nr�e����8Ȱ����7��`������ђ�f�F�x�h���;@k���ӳˀ�g�tӝ�$�׋K�3���HY�f�x����bB��q'P:˾��ɚ�B�{�22��	Q}O�h �Je�����7� ~�+����S��0��cw>6#c��&��t����#p^� I��E����̴�����:�Gu�g0@i^b��M]K��+6��S�eD-��d�ir�Ð���OO��� $Ќ��Y��
�~�6~aM*W�q��/I���x����,	㧼
C��l�y*�d[bs ��Y�W�-nU7K&�x�J���[���r�<�_��r�|��y!���?�?P
	㡏��(��6] H~M9��0�e
N�롔�^A.Ȟ،��7�W�c�|�;p��~K��Z-D���Hy����8+���0��0$_��Ε�^���>���3�y�g��?tR�w�A�ɴ`}��b����l6/>@�h���Ȯ�����b'���"����~"�3t�Ũ6��5/�y~��,<�){Ր,�� �E[����z��.�ó���ȡK':��%�^8:i?��_�J� 6��A�������.�E�ט��)�,����=V���qwy^��zǳ^H{�F���!��3��O�1`��O�,nA�'��ځ.U�����??+�L�]��Wׂ����]���ͳ����5�S4���7�>�+0�)ߘ=Wո#�l��~�O���Ћ�-_�k˿(�-�b&���ܨ����9u�}cቤ����kF��M�7�{��k�>�.Ac��J&V��e�X~ M�R=M!Kғ1�-�O4���Ĭ��ғ�F@���˦-0�Q���a�%K��Լ��%�C�GnF�~���N�XO�����m���nR���Zv���fQM��T�9%sr+�7E�ɁFy��nK���UF�f����.,]�8����[�ҿ�`�O�4�F/.��(�1P$���@RU�Ә�v�͸�V����x�\�ځ�gV�@���Qw�	`"L��{�X�����6Zmrm"�_�X�l�|/�����ҊҤ|���<�y?�F]�!0GJD/��f��k��Lݎ����T����
�`s�!U���m�ð�U�C�Q���1�';������Q���N�G�?�n�MbN�&�NhQ������O�gJ�"�\lE�"�F׏��x�j&�S�k\W�[�F5�7-]:��������/�^� l�	���n7e)�;��%^��|R�����~#����maY%��8�26P�*"w.ùe>ߟx��f_���S�C��öZf�L�����o����K���@�����FEre�P��{���>F����i�P]v�,�c=B2AF��cy8 4+�qJQ���8���r�2>���-�մ�p�LL���)_��0��JL��ys�%U�2�7;���S��Ca �Y�k=8�<�x�ZpS�`>?�unZ��m�)!��cQ��+��"mK�:��~z{Zx��l����F=j&��C�Ѩ���G��3��C�ZZb4��>ֈH�G*�X�ƌ.�ϯ� ��[z����W-��j�_ٝ}3�����n�[�N�f��T|�Q��~<���;k���/�q�puF1�X�}������g���7��LGr���ͳ74�N4"�s.t�e���h�-��I�� WdE8¦��#߀x�1�|�-���7�p��zѵ�1�ţ��fT�_+^��5�09�v�r6���͓r7���S}I�MSš���c��#�������Ƣ�����D�j�{��8��ױ95�a���C�t]�2[��4U��l_V���"H�~����8��q"���#�;�omD��6#����ו��Q�G^p&@T��O��7��)S�S�I-� ៶�«vC������wR��T�z
��wz�ux����B\񥔇�B�@�K�:�u/�5��霍�����:M��c��,���ç��JW��`m�۱���uz��I���-2�qu��{���)*��2�MV�}�ɵ ���>Q��G���QҚdQ\]E��ِE�͏8��|�p<J���������p��S)�<�U@�|�f%*��D,d� ��v0Y��x��f�tv��NMC:�u����� �L�T�\�(}��cc��D��b'�YK��X���w㸦�f�t,��S=�.b:��H�:���@��2a0���@rj��c�ʒ�/nC���7��,�T�%\ݼ%sW��|_����C�
^!�$���"\�8Z=_;Q�wų^�|�A�.�A	����C:��=@�w����7Qw���낯��ބj?����*;T��澼����J򹤣�h��ٺ������v�C˘���$�#w��_�Ѝ�a�a���5�e�������N���ڹm��Q/�r��3'��s�G�31Yr���3=vt ���(����jg�����d�e:�^kq�LE/��j;�(=�u�<3�AU���=�xv����$�͗-�?:G�G4֯?(r�6�Zyy;b	�^��i��U��)r�uس��{�G��R7�8���NՉ�q������}x�R<��!����RMR�)���]sW�O�Ҹd�:�eC}�I艭e��W�O�v�>rZИ�E���|b�h�e����C�?;��%�m �n�];UW&���4�:��3|�J�шS���O��Mb��ŕ��vT��O��U��&z�q��_'�߰�d
0�������W�I���� �EU$hDv���~�^7��e-���������,�/:\��_������Vŭ�p�2MT۾<�r}p�Br&��یOw-���yW#����D�-������j"��H~�� � 9a�g�\���z���&�+��TG��Qp�GY#v)+atq��EJ]�����%8�.��nt0��P�����j=j%���EM�v�	�p�~T���;mx�A_�bK��)�ܴ�xJp(�h�h�`%����B}b��J��^���X��ؿ�5�
�,�˓�&�R6��O�tVK��:�v�zwϹv�\�D^��ɼT��x���VpO�)\���;DM��R�sax�vm�R@���W�=tR�\2�A+�(��Np~�!�����d)�����}���}}U��i�PQ�?8�
%�.��ϯ�.s��.Xm��z{J\08�7��,P;+��c�u�zΊt�芛(�5n��{%�Zg_��w{���v�];�(��b��U2s k���A���o,�d����I�`y{L��̲3z^��=G��]n���ku��n[�1/�gq�#�<�Q���H�������is�|%���J�𧻓&S��VW�(�=�ch0�J�E���t�1���i�u)^���ˎ�j�M<�q�;���8����ʰ�ypר�G�c8�p��j�c��F�M2��.`���]��)��[�b��/�%��%������oBxjR��4�"G����(���2}��˼#���7t����Ƨ��>��j�g��6�t����C��iO�	�j��A�rl("��ǧ�;4|ʱ8��C��+7��VC�+�=K���&����0�_�<��@|��x�ۣ��}�v���x]�Q����L�=�<�
�����c�hx�r�3����Z�Ï�9�Qztl����v;7ݖC��O􇿨5G�ղ���57#'�ӡ�r������䮁MsR�rX@2��˸F`��bķt'Q뙔7��:��CԦ�,h��XTױ�A���,�3�l;��Sq����oӝ�!b9��� K�g�>�N�7Ӗލ�꒽mzA���^�!�e,���&����U��������/q�FC���1_���"M��@�`;�Q���3�����Z�z��^�y��s��}h�ߛ�!̬?��64qe"���`
�y����D��ს�.?�����ʙ'�����Q����Z�
����єs�B�Bf�����U0Q%q�c��H�]�ǎ��"M=U�;��8�N�0T/�~yP^����dy�]�b�]u�K��	w�YC�@�պ���}�oo�⦛ej�q�4�dI�>��3��E���E���4�1_7�aɃW՚�W_��l��6�4|ThfR:5مf��S<G�Q��j-|��!�<�z�5�C���7�O��A璽t��JH�T;q��X�FeR�7�g���6�L�m۶k��/A���f����c�	�k���E���	�>\�j��ѫ���\�6\	�z+tt*���6Z��~�h�y��E�Y[mwx_f�yD8>׸�q���\���bI��%b?�~��#xsG9x�|�\����`ڰ�����tH���ݏ���S�l��͢���t�0� Y�U��	<ε��UII��3���m�ZٰG�{�K�S�(�T^DH�����jA>��{'��)ܷ�=�g���!��4���o/"�䅡�}��^�A��m�wϏ�#3Q�^o������������U����D�Z��l���틓�iH�Q����O�I0���Ҽ{�vϥNoR�!��M����]�L)4~ռJ��CHn�&ʊ��"��,G�@wx�r�Z�/�6d;p�%~�+ZHC;�E�{gֲv�u�Rp��C���`#���8�w��ނ���"����g�2[�~꒿Y�FQ�����oR/�y��}�oJ�3(�zp����ߙh���5Y�ܦ��`A�)�-(#��h�����Y1�b_b!9D�U�j�O7N�C`�1�vz������7[�-2cTO��ֵX�/��ѵr�s����I��K��H�J/y�T��/�>�X�^E�(_�WȬՍ@vten}VX��w�ԼMk+]˜u���g�g�)O�$S>R`F�6�=NA���.�N�����Ҷ�׊�B��Ȇ:a���QJ�AuP��D���IR�1��Ui�,/�b�c�Ȩʧ�t2�`�V�1�J23�7�7OFT�WO�տ�KQ�io�˴�ͱ+�%>eiǆg��@�����Ǜc��d$y�.�>�XV5W񨸯N����ˆ��4%��zt������8d�0ЇɏK�l�~!1s��@F��|���Q����Mc��ލ�n���^�l����%�n�,z�S1�tB�aO�/c]?�U`]�:6Y����(��WP� {�o�Yn�ґ��
s����I?��9MfKSJ�A��vdC�Ŭb��ڜi����<v�f��=c����皀��.�0�n�#t��o��~��~~$xA�T/���AB�0�^��䡑X��w�ɲm?ɚ��)z����9�A�1��H������~mw�d��n�������"��a4ik۳��?{�\�4���c�����I*$�lB�Á��fw��y�mc��Ƹe�a����5	m<����}�YNI^�Z_�0���{^P>�n�ejd]<���]Gn���[\«�֢�&;V�Ov��~0r'�f�_�ވ|v��G�8f�uO9����3�2�T�n��a�Z�7[S���/�ѐ%��6�ѕ�H�c�u`͜<Q?�Jeq�
};�y7��D�g�m�}�V�m����ͪ��[��ǔ�����F��s�R�qsh�E$�5T�����j䭉K�K�����]�R7x����>���{X����ƥ��WR/_P~ˈaE�shm�[3���3�~�q*r(ֿ��9A��Ufw��L6�m�`d��)��+��?Z�R@�)�
�Bb��ʕ��9�W�w��^�"�i�O܍�U��v�0�$�^y�D)��̅wϝ'2��x;qJ"H���F�T����a��]����2� )����C�}���YI׽�]ܙ��ٵ�o��&E�7��{�>�.:s�yG���ܡW������سu�{���(f�p��.�Y��ǆ�Ų���vv8���Hp�'lhcGޚ����)��}p�6�QY��!���v38`�=����,W��!a��Jss5�N]��U1q����c����.01�O�I~5w��Z�G򳀈t�>8ރ��w06��[n�/����,�<������w��(�UV���O\��l$1�z-(����uj��/���*^`�����l���V|w8�NT]��(r�m������:�ED�rE�as�abm�b����q�N]�����s��_3-�1ݤ7ӥ�l{$���*���>�K����LKC|���?L������������7��a<���-?�<k��ų�TV@&!~�b�H\]��bu���vk��o.D%�;�P�����K��_;�w�<x9�/�B��Y� �s���|J�*p�8�3���k�qaZ]!�>`}���Wm�$��}���(-B��O~��T��/�)7w�>�H��o&�N�w����+ �d�(�i�gP�����$wŚ:�@�O�*�)�KԷcu�+�Y�&�!ʾ��|�`\U1��VGV�֦��3�r�\\�wX�n=3M�%������.�ݰ��1�������"�R������H�6���vj��ê3���%�6/u�;B�����nT{j{�1���u��|�%+��W���6K��M��2��$H7^)��2=E�]h�wN���~	�����4����)5;�zʬ���چkv[��_F�n����=(D,|y {PGt^�G�j2��=J�QQ�\��bq�C`��<���V��a�B�أ�CS�b��,/g����,����6m4��-kF}�����.�u��o��vn���]S��Z���[u��d�&H�ek%�)�CB�|4�V1����cO��N]�����lUbv>X���l}���Y-e���6���?	T���)��?������/���z�n������M��A�+��^q�dH����2{�66aMOv���Mr�؁�.P��k)E5�iS��3��	C;���T���>�5���Kw{��[�����th��+�����c���m-oĒ����3���t�������O�E���[?1�8غ@TL��� Q�w�[��6z��pd'g4�� Y$]�M�1���.���׍�\狷E2d�>:i�tA�|��y�X��c6W�rh fn�����=.�zN��˺��s�����'b�5�܇3#��\�EF[���A��_(�s�ۚ"�<�"{74�W��4 Q�b�^�:q2���y�W��R��v+�)Z?8w�s�ߩ�a/�X�$2\~�B�ӜDY��^|2���&�]���Ii���4�B �C��O�e�#��ڄ�;�R𺙻U�%$�:�y';�c��MwW"n�O���v��"*�d�JO|���I	5���������������n����I�%�:�â���H�N����9���H�;�t5c��hNUc�K8�pEyy�}G�����c� �S�ysfr]K�.��{�ۊ��t�܏����{
����(��Ӆ�M����E�Evi��
Eq��Q�
����a�p�=�u2ΉD���rt����t�߯$[?���r����R9O`����p����!3���b��$2Rʖ�c��ϻhP ���I3m�'��v'G�v���,��CO��/�B���='�k��:��ܫ�M��ȹ⚸�ʧ0��A\x�l��~�ǘ�[��/��=xdOP�I�JRvW̷��מ�����A�~��ܫ�HW�텭����+v8#�L,>-=��\��2�M3(O2%���ʊ<%G���T��g�s|0�K[���t��#b�"'�m�bme��(~�P%8��1��#8J��q�Bq�`�@8����_'�F�Mw��c�˓փ��7ONHY���^��_��d�=.��I_CTEn������P|L;\�_�Y-�D�*��H��IW��J������O���Yc?�sBc���=oB�/%��i�5/0�]��n
�V��d�>�`�=�4k���ܻNHS)�r��}7�/�O�9_y�,�*�"�-4�Tix(0��3WG�-��� �̝��cj��'����Ձҭ���=���H���!���O.��U�%�B&���u��Qy�l֏����3��`K���{z��[�(]m� ��VX~��TY���kE�d��cu��*���y!En�ڷ	��3�k��R�}�Q}��Lιz����g�dB��Џ��M����'<}�Ebn}8~1��M�>-ɯ:���㳰fY8d�Չ`��A8��vc�?��Z?��U�lZ��Ӣ�3߼���I4��n����Y���ƛ55�Ǔl�̡�=��_����Wx��M�gW{k ��֙Y-������H�CW�{�I{�jRհU�8�{��L0�ق_:Rީ1&��I��1\�����8h��e�IU � �>�r.��]�Ի�����M�_)"�A�-��p�\����^�����H_j��:�H�"��F#�B�w�y����|
aW��zb��ibF+�����ݦs?�:
fM�2�4S51��׊��͸aN��1�@��~��b���T��9�;�8�U�φa����r�J��I]�EU��������s� Om:��	�
��E���+B66_��X̚^TeX�r�=*�\�� �@6���fQv�|dm�JW'�L?[}^�^�1�a 2kYUܞq?���ɹj��WH�;�� ~��ݤ�?�EB*�0����ٍ���_�%�s�'�y�Ea�%�݁�8����繘���/XhY0�.��xg=�e3��.�&p3Z�����	�Ў��z��\xN��e�|��_�$-%y�}���@1��?5ϑ+3�r}虍٢��G�Ua�#sϏ��;�w��O�UkϻW�_�)� "a��dY�h�з����C@��ςdW:�T��[�m��Ϩ���p#���ů;�Zm%�j��4���B�6�C��3`F��e�]��xƩ..ʙs��6?΂������)�U�W�[N����M���wk�ŏ��ǂ�B��`����]����'�V��\ТyG�P��qT�sX$���!�+�%A@�.����S%�2M�P88��f��������^}8^�����{-/i*2�#Zt!�mM\j`Q�:3J=����:|1�u��Ud���i�/Վ���M����#Up>�g��_��X'E�:��HcNM���+��d�*���k+�p��{ ~wE���"/� ��lh�����j1���E)��>�NJiwk2�����\�G�D��c{��B���N9��T��?�(�;�{EݶyҹH�1�L�:��ZJ8����������A��1��鷂7�gȂ4@���	уB'��(l�/�R1��=��]c�û��!��&nC�G��Y�(�M��镇����;V�"�e1ɤ��J�V��0s�nNw@9�mUX�=0%�Xꤛ�Zv��^9jA�Q�d��g����d��^� ��I���w>ͪ"���ى����[9���4��$� ڬAm<�jj���G���@O�o�W]�bK`���������8�0��-�<B�_&èl���r|W�asM08��8�	����X���pxs����?�♱�,W��5%�Fu�����=�~�+�zf�n�m֊�2���<�9�Mr�r���"@��"gX�Z굵LHɿ�g;�u���.�%��o�7e�-WVnlt+�]YM;tB�����'�F�N���Ԛ3��`[\��le̻3`����V9�<��afH��jC%�6�Ćr#}��4�Xڄ|�r�ړS�� D� �K�ԣ��["��Q�O��Vj�z��9|Aet/�?r����p�:ƕ�6I4@�c?�{P�"�:EX��_.O\|�^1�=�Q����1�ۅ("���)���9�]��	� ��4�O�f�b������
'2�٢��兏 	h���H�*��R%����
�R����g�Ѿ�eҋS@T)j�I^jq	�J�g/�����=R_�Tmc<��!�-������[O`ޫ	d;�]ͦ��/������Q�z֑P�M)h{A�-KL4��1t�JE�q_���`�����G��$��>���3'��j+�2�s�x%0�N�K<��U7�t?h��Itu&�A��m�`��&�Y�k��1R�ɑ�9�*��+�1]i�=�y��6��0�Q�u["�c�g����E�
k�`K���7���5O`�@ׅ�"�,�Xf�NB6����9g�Ir��@���G����~��+���k�iFHR��Ѯ]�j2��{�7�6�����	���h]>?�>�[��E7���9ͥ�=�3�	��d�'�x��7���,�Vj1黨�Zږu"o��6�{^a�����:��d>�A{��0�R����m�L���΄C�^g��p]G&�٩�&/���b<���o�f[:ww[�nX�E��.����y�bN�0�+:5��M7h 1�)g�)�מ�>���%��۵͑�A��`XcD�Pg�����%�r��0��[��';\��M�z|r�&�D:Ģ�t�:�)�Et.���/i��sq��
�zb��"��l�0@o�Ɗ�X���a""���F$���2?)�A�))��`�`2��T����l(�A�:~�b<q�&v�mw�a�D��W��Cٟ�+\,��3�ٷ��b3�fFy��ݢyI2g,e�V�� ;�>♓R\��Y�9̦�_G���Mz8 L��GR��ݤ�H�O���Mi����8�<mY���)t�S���C� ��_v��ds�0��g�)֎�A��"�.M��Q&�	%�A��q��Z�=A������A��V?�7��=�=u��yQ+�8k|_�FP+�.3-q^�\����to�O��� ���H��'O���G������Y�Ä��h�6GX��Yd�ց���,�M�� �*M���Iv.�ة.��nt���KR�F&��^:�O9<��A�'4@H���qx>x�Y�8�!�����[~9|<��d+�؆�YiR�UC��J�v2���(���~�oG�7=�\�i�+�js��w�R����"��$�5bZD����H�u���~O�h]`���"C����]�+�����:�C=+P���H�`���Q�Ӟ�E/���רj������I�Ծo6�-o���(ɿ�"����2@tƓ�w*)ML4 �H��߱�?�X|�������#`s�z?�2vp�
i�\��,�+R���x� �h��h譺���';�ar�����B{����E�Az$�R�N�ٴ&r"�f�ŋ����t����"Ɖ�o�5Y��K�[�u��i>�_%]+�������D)L<��t��@�EAn�_&��d�-��?����o�z��O\컎�u@-ԘQ�2�B�̩t�G��\Ҏ�Y}��c����q5�<#�Q�� �5�6�@%�cB�a=%�ɍ0z�TK��7=�oXT�ٻ:�fX��pk�?���.�^	Z�qMi�^#/�-����i��?j�Db�s����B���v�-��0q�UW������@��</ꋑv �1��� �&�P��.�D 0c�e��t���Gҝ�l����R���tQ�����<��F!TeѢy��ڼ�vx��I��k�~���׸0��Č��y
ˈ�Y*m α��_D#ڭ���ꢕ��^D�6^3Z����EiuH
�1p�h�œ��;���\��i�����r����h������).ӷ��/*�<����O�,�e��le7�6{�����[����	!�,Q���2��}ɾg�;��f��}~�<�����}�����z_�u��y�W_(<7�Cn(1yH�%п�YHFvܩrf`��Ή��MQ�Qi�Y>�|hz�(���d��H�ÙLE7����e�*�a�q6��5�e�����ߍVb^*�&����_���Q��i?8ojOM� ���^f<}KTy���t^ؿ�o��B�1�U��8�~��k���~�疕�؄��W1��,�G�0�/�Ց˕����h��-��1�m]��&'ÅKn��P���1�H����R��g�y��G�>0w�V���L�*m��)A�\?H�c�����a�k�p�i����η�pz����l������G�{�j�b�W�G�� "/!�񓟄ю��?�=!��
b6a�f{������>�d�8�ƒ����eT?6����K3!�Et�{�$��k1Y)�qC� ��m��W��ƨ3E%��a����bTo�L�%�m����tX��]2���R�m�Ae�{��ڗ|��g;ӣ�֜ړ��u2z*D���f�\%���b��1+��r���k��{Wz<���9Z���t��>g溏->�p��?G���h���	�/7��%뤌���)O���Ѡ�N��c�\���B� c/�����C~̛i(�W�䑥/^�f\C�08)A�J�[\�fLۖ�q�Ǹ�؞iq0�w��c�O��ɏs��GnL}���"���߿�G
�ݽ�$��x�i%/17�9��50PV��Y��r���=���Κ,���P1��e�֌K��{��J�c����=4ư�u�.&�����S������.��n�[b����a�T!��T��w)���y�N��8b��efH��s��g��	�A���Η����^Ѷ���oT���y��T(��ݑ&��%�{KC��1c�=ԧ�F��FW��R�{S8h��ؾO�жW�����zۭ!�����(���s�u�:��X�'���iS�j&a"�&6��k�p�>�]9׳eX������%��Zg[��1' /��Lp��cC%�[lIU�Z�����"��=J��|�߮��g�8+Ւ�[�U4�������:�n0��N����S˺09���R^�+:��b��S��؆�Y�gpz����o/���~=�_��`>�)Rq��� ��@q�=f1V�.su�H�O�+Vȸd��%5����]��2���E$���Ku���:�
��'|h�q;���e�Κ�����z�}sj�v����l�uҙ�n�;LY����-e,jiL�:�������W�����?1m�q����9�?���W�	+F}��(�lE8�ޠ�Д��9�q�@�	 �I{�����+�����z]M>�_
�w?���Y�;�����.$�S��t���b|�"',�!��P�2g����.cW��1G��,�M��UN��3=��P���$����Y�� $vM�pC�*T�x��ӝ������DB�ʐ]ٚ�M�����������(��c�T��Z�>с%CY�x�e��r�6���9��f�0?:5���[XOѐ����������t�%����"�!L���s�I=�����l�D��\�-����,�;����?�('�l
|�Xv��B�G�?��M�f=�2��r�}��a'��{|zU�s����:DP�1y({�5��|[��P��������� �Vz:��OuI�TE��]�b3;��W�5Z[EJv��8Jc�X�ɯ�~�V>ւ��$oo�m�ڿ��a:Z�s��SQ8`�h�q|XʂT)vp��y�;q4u�L����؉��a̟�2=V���SkH�"�y���i�כ���4Gf_�|�!��@�y� f��1�)�w
Yٌy��!@����,�� `z	B���L��9�G��f_;��t�-f}7�ޝy������ Y�҄���ϊ�}�[�)�;���IBg
�.���zO������8"
��KF�������K�b�����]��,�f�Br"���J�
���>}H�L���b�ΨA�S��A�A���`7��ۇS_j}o�u9��Y]�mG��~�B��^삲,!�3ya��GzQ�A.7���U��O�w��B��S]%�<�b��WqV�)s�4h��:c�t��ұԫf�bsm:���S`k�s{�Rp�T����aF|:�Z�h�0�+�|�J/(��#���L���B�Ӫ�\�-[QF���y�p���U7��U���[��&_������FI�M�y�k�d���<X{����.�����R'�z�2���ɏ7����M�8��
�?}>'z�x�*c�X�8�[D�P?A2���);�e�y�������M�IGҤ
O .��1�����ⱂe���R�~ʴ�>O�=���d -�;ֺ��ѥYӋN ��Ć��\o,�:T�D�|^��zIHJ�sPŶrB`Cj��<7�v�$��}=��rT{�*"EB<�/K��-z����Xm3���B0ٮ��օ�;�\Fr���kՐj��E��P-�"���P0�i�=���`����Ps�#��f���oxH�߿o�7I�.HX�{���*��Dά
ݗ�JM�Y jr��ty��$F�!dCz6�]�1�X�څ�9�M{��o�o� =\c�,�u�..X���8���.��/�fv�ݵ�M��8O z����XvC���+��#ۖ�2(��@r�iB\0�-v���z�ƾO>��Ѳ�pY� �{a�Bo� \O]�K��Q���e�o��:�Z;�֊���+�~���� �����rN�H�n"x��׌�̻�f^y��c�[�v��)��SPj(�BE���,H/�.vL��� ΋���.h�ڥy�8��1�_��X��{Z������)��)���5�O���͏`�f�CY�n�"D�(�YY,��$�n��+���(�e�&}}��H����f��IJ�=Q��*S6�"���z8{��㠱���ك��Q�ȝZ%���tʽK6㵕�
W����M牄�j?c]>�*mN�+�4L4k/u
�~RlEm=��Sv�%G����t��>���G�yxi����vsHn�r�cc����?����;F�+�諚a��P�[K��U/��H%��Ÿޛ�S�Ry)!6�����jv�ϲi����f�Yc�N��|����y��`��u����ұ U�Z��j�@�1�昭������Sq֚�y|��"*���SiF1��V�U�?ў;���(�� d=��ݞ�SҟSDs�\g��vbӟRq^��e]�oκ�貽U�ndk�ׂ�P��o7&�?�p4Z��S;��񡷋���^}R�
�5-�T�������)6�R�iZ����&���ی�"�!_�Ez˃��?/���s��v�,�=߂�Z]/0��?�և����L,����b�~�M�F���+��n�r� b�(z��P�0���2q2�\�~4���j"__�OE��a�ܟ�sxj���H:�!@��az�1(5��S*~�ի�}�p��P�+,Ѭ*7��\���Re���Rs&\�^tw�� �q��Q8�a����1������8��T����P�I�8t�J+\i?���]zߝ�Ⱥ��0���#F$p��������ha�4�#�B��b�����%�s6]o������ �g!\�����H�l��ԛ�M��IX���d����*�_G��c6����^*�ң"��Ӑ��?�^k­�|u��\�J�K�aB�������|�=�OD�j-G�)���z���?���ϣ�a��z��S�r�)\2�2�����E�Ml /��´��b)�f^�^>/-��d����zKp�4i#�⭆�4�%�qc�LҚ1�%yʜ�E�*F��P�LJ�im�_����c��&�G̅?�ҳ�ظ��%� l��0�%�d�P�~�ø��pyd�PGa�I��'��?�.�����c96�^ �[�@��I�居v�'OC<��l�R��9T^$�	�ާI'��Ķ֘tI�Hb͊�Z����'����� ��c%� #�zWlZ���;M5&���j�
��p>�+ܜr��Kv�g�A^9����snP�ۚR�:�yf�Lޓ��M�}>�c��&,���e��|Ppf"�B�Vʴ�Y]Qҍ��8\��\���#����^���wO���덾V���-���Y��ݼ��l<��n8��IfJ'���X+r�-�~��@���@��5}4l�q�@>Ȓ�6����?�����#�>��sO ��8���ߙ� �s�SoO �\�� �1�T�T)��qg9�t�Z�H�F}
s�v����t���Ǐ=��YH	��&F$��->��`-?��ӑ��N-����[�T/�=�~�C�XK4k�E���A�ZЅ�k<K3\1�"|}�S8�����^!���v����$�e~��ϧ�a�o�h�;�jY���8a�Nߩ6���N��,��F:��$+��� �'��W��W\�����煃nk[���D�=�L�]ҫ�S�8<ylJ"�0GjF=ǃ�Y�3O ��i4�-�c�3^������Y����(s��<�I��h�I�M�e�p0����	��$=��7��+4o�e.�/I�[�whT�����Z�&���<]�	�5r{�b�����k������}2z|�][�Y��Y���P{#��Y���k����])n{�Y ��Gg�.�N|�)��,Md|��qZŪ��c��B��Q��۔Jc����y��~m9cr-L�Oag���Q���T��F�Qz	�jZR]�j�����]�1J���=Yd'q.�C�^P5���Armh8@��,؋�=m0��Y޳��о�$��n���"�}�d��D��5�9����T��b�ٴ֌vM�"q�̳e�ڈ_#JuzY��Uj�K�)[rq������lz�.��g�R�(�SZ���ey�]�.���F�GP���B{����^Kvr�0���ZMou?��U�����H��X��w��?���]4R��.G$��Ձr��rj@�$ir/�0�� e��ra3[l���o��A`f�����m,:����_�R���n�%~��3AFT����~wI��̤�M?�b��i�K��~����Ȁ]d%1�� r��L��r���o�����Kԩ/�N]M-���3BK��a�ҽK�������O���q��?���z�QRuX�� #B��o�R8]���eX��[~0K�=io�Ob¶�ǏT�<H�(+�'�{N|v}�~v���A�o�b�h剦�����v	��g�sŴ���Dꈍ��BI?=}76}J����q��/I7ߪ�v��2\�:	��`J�!l�������t����ئ=5y���������U��dۿ�$E�R��p;uR\�V���!�y�-�)u���9��3�����x�N�x��(���,�WGl��DY��i�F� Y�KޫG�:?|G?*�^r�'+e�>%� �/ ;�B' {EC:�A�:��L~E����/�ͫ�#8�S��P�8%�`Y�؆�ӡx����TC�MG����s���^�-j_�����)�^��lsf\���p' ��?��FD�T��J�AX洏���@E:�s>3�m���5@�g��t�����7T��̓���M;�m�ut�+#����D�{��U��qJ}E�q:�� *+�|e��y�1b�����9��e��)a����5Y���� >'r��%�Q�p�(�I���kS�$���"�v�������b�	�q%��sܶ�?L��7��D��	P�Σ�&k"��J��!���Ȍ�f���� �4�?'V���񁧆*�Ր�w��1�-�BPgص<�O�{S,[ �<z/<�����GHb�1�N��r�FOCɚ^���=�����sA�����p�惝������Ѥo�w��,'�j5�c�'���J����R�7��(�k�E"�0��I,��,��������x�>B�?�ʢɔJ�:�v-E����v�48��P�:j=? P��s�x����I�m;^���P���E�lw)h�<�����#pq�(�c����ǅ̚g��(r=��f�q�M��I��(��M/�rN�iWY��:��� �o�2��&`1�3s*�ZTVNޫ�P^Q;q3o~na�/���T���>Qyζ@�F�.��9��B!̹��#��0��G�+���/�M'7M�E����ۡ	�tn����9�Ӿ��Zh��C,��ٜ�F3Jױ^�4}i��X�����Ucrx5w�,�s�,�o�6kÇ:O <��)K�(��n��F ��=�Y�t�lõڂh����,�U����3����P��q��~�P
y����;��D�	����5��~a׶#��H��{��M��y��UU��Wd:�����:�`���1�c6E��Ik#A_� �lw��lt\�E_�=��Kiiw~w(���x�x�a���_J-�rPq
I���7��4il�$k� �b�r��	`KiG�ާ�?�W�� F��P� �_�/�B�:��S̬;�^[T&�}`�6i��iH����9M���wiR(� ^��{Z�}���D�����#@[7�E�z�kC�7!b	v��9�Q�d'*���_ ��k��'�b\��Ӧ~�?���_A����Aؑ�:)�SX�b��Յ��3sv���|�7;�Ѽv�/N�\K_F�R|q�2��jTmo5����~��;�Rm�:2��P���64��
T�j�pH�U�j��m����fes�S�Kx��A*��C����L�"� ��N��_-�+�Sk��]X�\������+{x��\��lۜznD���Nc#�LE�s�� �S�R�E�7ʭ֝��� | +Eb�m�!�����0-<�QPr<¶S��"u%x-�9݅Lh�@���p�yb��g樚��R�����8LrJh��6�E�K� �q��8���ah�B�}�.'��ʏ,Hcdu�@��Y�xI�����M%����Agm��?]/���8߇MK�� �!�D㥩h���ϸ>�oP5�|O�2m�DV�t|~��'�U��*��\Pȝ#�ҩ����..�"���w�-�'�^�z�Y��������Y�\f.�w��'�lh��T�Ѽ���(��N������g_�BU'��}�!?����18��Z��Q���%$ۍ��|}�3��_�ϙ����L�� (X�el)��5�2��[A���&�����>��<�r���2%A�~KR���M�*k��{�O9x�P!�2� P��4>���g��Ù3z�:�.Ϯ�O�����qNy-���4s�h5����ׇ� ��-R��Z	���'��w���N���x+�q>����g��Uht0�q[�P�r�÷9-#��[��N=s�|�>{�|J��j�R�I����L��F�!��	eꥈ;��LA�w�r�̎x�v�qr!����Q:����+0f_<OT��Nm5�U���%���H�<"�&�3\P},��-��!�Ec�;$�^*�i�3�l-6�u׾}dU?� F�yZ��jk�0Z?�ZZg/����9d�{	7�Y7������p!���w:�=kR--�&��{i�^N�C
<߿�cp�D��r��_N�a+&}[dpm�w�D`�=E�p��\���A�]=`2N )�OW�6}��y���oV������6�����%�r9���犭Z�w�+O��!�m��ҼN &P�׌R�i��i��6�*x������L��~e^����ذy 6U�-��������Q�8��W�I���3վ�p�/'�D���2-� ���#Sa�o0ΤE��s�1,����ǖ=�Hd(p�v�+��cH�ġ�:����z��x�χ���#r��%OWE�	�]�S�n@3���6oxv�Hv��2$}Hah"�c��/]���C���Z����~�w�u����^��}���RXB�C�5߰���o��>����a`����w����mfe��Y�"��&�ݛg�S�����Z�U+�b��b����
������ّ��V*�Z�z8��m���1���VC)�� ��'[:��2s���I>�9
YS���k�f�H�5E$�N ��l��͸B�P�-a����O�n�%n{�O��������+U�/��VOB[E2Q��\����Y�o���&��K���-g)F@�{0�[�rT�v�0�Q�Xҧ�����TaP��*���H�[�⨁k�;���-�ζ�z@AYr�B6�ƅ��>�+����#�"
�F�?�Y
��j�,�9T�{�˧�ן��.V�N �^ȗ;ӱc환�/ڝǁ��+�����^&)��ʅ�٥J�]|���p��S��7�hL��+A���%h��?7�޵�1 ���e7��į�yx�ԌةO$)>$�Eނ�6�N��ǩ{mg�'���w;[�
,��o�P��QS��ݎ�W,�|Po�:[N�0r���H�Cȑ3�_~HE�d�~��	�*�8 ,��z�{<U���ԙ��"�&p�V��N�����
�:���H6����,�C��4c7v`�[�������B�O��ڡ�N6[� wN�`��0�1�q2Z����t�༊yK�?:���t|(~�$���ѩ�3}i��~������E��H�lX��Ll<�N2`�G�窝Ul�!�����0	&��
1��x�z�A���Cg�S1m������X/Ō��[j�'�Q4{�m�T;����hi�V[�s )���ܩ��5���?x�5x�ր�t��o�u�ѩ�j��d�	@��݀.F޲״7nN����y��B��B�P�D���xp<5g�|����ˢ��j��N^�=�QC����<��+�',��y��4DEq�g®�r������]/ۖ͝a���R�(��D{k%�}��y���j$�GΟ�E�$����s����L�.��Qï��H�G:�`?M��;�~vɩBO錞���K������W��l�䃴�M�L���,cm�'�����s���1JS' �!1
���xH0+2��Aa6k/�yUt���x�2R*I�]H�עb��;��MT��Dc|�t�RW�|��?�T��|�&]	sB}�Wz2wW/؊ۙk�V
��!폞m��}�r�S]���(ZyYڲj��$�+z|�׉����c�P��ov,m�?��@�9��#池@I�vZr��RKwx��^�}����&H��h%>Z�H����nv\$^l~ޤ��e�l�D�n%�凔�U@�D��@|�����9�Op3!1g9A�B��XW�`��I­�i�F�![�5�������N(�V˽׌�W�Ȼv4u䓴�7DGٳ���
��M��*JcO�+�/�!}2I�g��68Y�� �Q��j�p�ɯt��˻�Ϭ�g)�WY�4�7OӣG�\�+�(�<r`�-2�%�Y�U!+u�g"r�'U�G�M�I�� h�!�hv�Q�L�ɣ�<�ٳ1�_�Lשׂ9*��\&����z�/\����g��i�]��z��*<�`Uy�o.;�d���%��p�.��[Ί�8����~a���� ǟ[�V#�;bk��V\�rMSXՁm��{� ���w��G.��4d;'�� ڽ�� ĭ��������,�P�� >�� �^'�`�U׻�����S�������q_���R�tC�H*�FՀ,�R("n�u���M>xa{&�b�?����6�I�f�i�v����:�D�vk�
�;�n�g��dP�5�J�n���v�T�����A��ڋi��$l��;��b�����ǭ�a?)Ϯ)���^h��m�6�/~�s5�Ԯ�3V(�k٠�>�����|�"wgMz�\I�PE����i�)�������ۧ Pw�K�%_�~Q�?�auts�M�u�͎��$�YX:�k�7Å�)��=���=S*^�x���w���z:�m�5��&q'Re�j}�����[�cHn�bHU��K���U(f��֥�30hWq�B.(e��G�����RΎ��w�
�6-���J�i��"��,��ݛ�;�h�����})� �����'bރ��Ѕv�d3rP1���Jt����]��9�j��р�!�X%�� ⼬Faf�������S�_f���Ew�V�ª.��Ĥ���\a]�.RB��l�'�s�U ��\�\����9����h�cLc��?�������8�7q�%�ҲS7H�������O��a;��!�P��QT2��Z�㙡Lm,RKפbp��!��Ǘ���P4���#B���T3N1��GM�O����=i���	��w.��}2�[�즕�`�<Y�z&�Z��-��hRb��5]�&��Q��/�*�|dU(ݽs��bopw�}A����z�%N~�Ϲ��
Ǒ&u�f���4�<��~���6����?9��C���d���ʕKvE\S≱2���(#w���|S���� �e$��g�4�WW��<`)<��?O)�I�S�.U���Ӳꏟ�� \,d*`ߓ��%>��Y�����Q��;�0dgq���9;MqoB��
g��t'ʩ}[��o�	-�X݌UϹ>�Q�]��W|-[�w�?R�@���?Ye�}�ǃ�Nu�b�V+ |��������へ>.�:��P$h����Y�u�/�Kҝ�fx�hy��&�%��F%�!�4�|�W.����I;1d�������\����
D�8�x��-nq�:bW�Y9����|���!���4�Qi�'�����En].i�H}��d0ɀ��J�\lg�����.{��0�yH��	�wM���D�\���Gy�]�zR�x,��`���{|s�D�X*Y�b�J@W���]5��G���$����*ō��T+�u߾XxS#^q��HFL��o�"��G��iM��?
��/���G*���?��φH�-�O[���%K(���t�2 o)^�!��)D����<����"���д6ΘHn�V
�)�E��5@���vg�`.�!�쳫�L݌��Q�	�Ti�Z���i�'����g���J|����o��v�����d=��dLl'B�����31�k�Rz�RXHN%Ȅo���2�v���u8ϙ�ep����8qJ!T���n������'�~��7�\�E��zh�.�v�����7�c�����.���{Fʏ01Y�O5v�:��`d'���!���D�}�B	`�=�����s�o�R�ς���i���a3�!��=�KMk�9�ڞ��nޙ[�V���\@D�Mm"ȉ9��[u��ʜ�m�����S���� ��,�'0e� N�#u�&���M�݅��r^
�z��m�j�U�Ȁ[F��6�-���#�����=�;�egv�َ 9�(�E'�Ȯ2!�r�6u��G���uXφX�@�.�"@�8mꪘ����hZ����1(Bm��/��D�#wO��h1q��|����mS�C?�^�8�'|���������˩Y߬��W�sf-NӠ8��(t'����=��t�g���`/ĳ�W(������d�%|��5EѳX�>�ݏ����7��x���Lz��=u�NB��7���(	��>�����%^ǞI@:ҙ�V]иtC��*�<6-���W��@���S������6�éeUI����~X.�=�u���+��6��5V�wЗ���zt��E��CLNϪ�u�1��D�>�q�G�pWO��c8�¿+ŉpH�<m�h<i[k��#���~İ7ѭ=��Y8O�Lo FUo������|r�E_ʻ���RvH�����2ӤI;%�yۂ~����޸���?���G��Q�V�vn�ʞ��"y8���\lrL'��~lu�r�ysH�	��_h���8~�|Y1.��ۂO�v+���~���6���X���� �a����1�����>�҆�M��~�����{�R�ߋDN�b����u�/�~� ���)+U��2��sG�]�����f2-pv��	d�Cňq�����J�e&��k�k�0X�
�'@��g&Z�Ql[�Y�I�S��E�硢Ou��A�?�F�&z�z�=<��W��ǒ����֢�Ա]����}L��&�pf�4U܅��P[�d��g���Enw�ag��:@8\�ٝa�2U�$��c�-���>�!�O ��ow0�k|{҄,:b���̡��㟅ɹLY���6����ݱ�l�98��֍۶��ޡ���{�o�c�ŊqU��ȗ�4�H ���)�w'@�[j���Z�z_�C����*h���K���o���8�8�.E����_�.] ���/S���G��@WA:æZ+ľ�z�����ZU��q�&�'�.+�]aP���Z�xbn<ӆ1��¿��ֶ���/�
�wG-�8�y�_��<�52H'/�9�s�-�k�d���� 1B�:]pV�@;�qq��[����8tl��IMT7���
��ͯ�9�RA�N-�^��\׏��TU\��9ִsc*�Ƀ�Y��\$w�&#��E��)�����<���o$���;d���W��r��Ad��iӛ�Ǯ��L^:b�@܍��zQ���r��ߎ	5�,���������ҳZx�7����3
/�9��)z���m�h�F�km*c���X���b�L,q`A#���"�p���-��-�u<E�Iz���+XH����q�o����M})����`��
������Br�׉��)�t������R�Y�=���'��RA9AɆ:.����1�1�)�mr�oQ�v�{�y"�xI[�=��͖P
�J��83�d5�vM�.�����]��3����I�R�bt��	��z|�<˓�QB�y��ºs�{E��^&��D`�2�#��P%�g����T2��F�ѧ���p���6o��¥֢�^T	��#
/�~!L��X�g�����b�1;C��^��?��~��F�]���C����$��R�u�����XU���ډ��!�F��*��1/�'
�̚�w��L�Z?�=��K�E�0[�D�L1Xk�w��"�#6G�~�z�;�h��#>?�ݳc����[m� �((�����������η�o��*ǿh-�遰�1x)!����������ճ���|�?%�ἧ9���q��������y����7oEy�	�:J;������ UdE&OH�S��;h�@e�W�,���'S��i'Й0gA�v~w翹��Y�U����	�D���߻�p�&//�
����N��o�2���r�f��H�$4�"�MJ��\s��)#t%�st9{�m��.%�	�������	�cpS�S(����@�
5+N�#2Yѹ�Ԧ���Z�C��:�p�~��}O΁�Յ]��ἇ�U��ym��vMD�k�P��-�����3 �j�>w��i�
�G��2��G�s���^��[��NL��b��U�)�	0Ga����͆��K�g��gNb]�(�$V�M�Bf.sE  	R!���b�ɟI0�϶x�q���;�����`#������F�ʄ�p|e��m	V:g��ߥ����~��s= sh5�Ec����O[�}J�d˦���'� |0,�K�5�(�r���V�`(h�؛�����K΋K	���Fr�Z�g�c!I�H+�O����:�M/�	*[���78=�v��ͱ�q��"_]1�W�z��>�Q\�k�8D2��Y���[�J�Zt�>V1��phRS���5�s��n���xE:Srw�u�����vTt�<U���p���w�~^�ha'�s�����賛�,'�J}ߜ�"y�R:��>L)��w�#w=�_
��u
R�C_���f�ڍ��������Zb�ی�v�z�\	�'&����x_>�l���M�jp���!_�$use��ϼ��O_~D�Xѻ�x���.h�"�� 6���pE�}�.+�m�N��D2NE��2j0�_�
��^R�\W�q��M9"u>&��Aǃn��j��xm��r�/�� \(���:k>�ͬ��:�U�<[�&~3��`z�G<v���fE|�A�1�������;�W2�i�ԑ���f;�͝��۪.�0ᓤħ��.̴3��Q���5�{/O�-��r�l���P���0����/4I���=CGe�!6u��O��!���4I�8��F�JL�������X~G5��ߡ3;]77��AD7H�� |����\�9r�~0>��0ѳ��+��T�H���3��$<�����}4�*]�c��Z ��y�L��}%�t���b�b׻l9
�	��@���b�}��Ւ-����:��\���C'%�� u�\�<����;�7[r���N���}
���V��h�"��wD�i�$�."-��+c��.Uu��w����Q�w�s�������d�J�b��	l�^�~e�� �m��]�m��Pe�`@��|���ٜ,b!��-C&?�X�5��w�����û���dX�[W�d_s���]a^Xňe��	�U䵊 ��� j uF���V@��5h���:6?��g'=˞���n��`�9��dcM����}�`�jҥjm.�_���A��@HF�ޒ���Q0k�oyS/��R�h9������j��t��)�.w�H/m�0a	qx(��z��������?��N�z� h���88��阴'i���a�	��˷h�G�co���cKjP��r�}�D|S�c��]�E��9�5��N���	��� Wɟ bT��=�쌿Rl����Wu/U�kX�+k�n4��yk�$��:�M�_��G���<�"
`�ɐ�zҵ����Ô`yM����2]��[��/>Q��C�p���i��Sݓ�a���(h�I��5M!� :[߶��H{`�b0$����r���f��a�s,�?tp����s�Zb����EqK�;\���������������L��9t?t�� m���[��)��]HTg�%Y^ש��6#&�$��"���y6Q�Hj�E�5� O l��x;��w�g*�/��
4\�s�8���D�50k`v�u��(���:�O�7Kw�������%��Qv��R�4�>��q�qR����V^Юܨ��� l�2�y ڲ-*�=p�ȽMOo�h��@t��Y8��+�B� ����k|�d�a�����2�U�mNi�V�w�}�J;�кl�DY: Lx�ص���.��睢��y����gR,͜B%F�es�Rg&M���k��֟����;��ZɖLE�+�b�|{-��W��Ӡ��Z�����-jD�(���)�*U��i��#�PI9֖V�PM�AQ׈ߣ�����#�jSW;,qU:f���l�YnM0+c��N��_i�Q�Uʝ�������[��&���콤��7�?�M�luj]������^ɡ|׽В�smF?���FQ�k���7�ʋ؇��C�O������B2�nzp5mR�j�/��0Ba�Y��/O��=�P����_Wtz];�o;Х��	�g3�<0�2;z7��]R��;�XIZ��J,Ɖ۞�9��P����u��*F�i����b�g�J(qXp[18,ӿ6��6����V��'��T.����v�Kr��<��gV�i���$Ё>7��ha����{����^���:�aX��+Ēm����.4\d�C�+�Tj�s���������h��M�J\���h�뛟Ӫ9F������s�r��UV��>�<%���,'6l�ݶ���Z�I9;�k��!ݟeE]z:ǟ����Ս�(ˡ��V�Ǫ���qBO����fƤ�O�:� b13��8,*������"�fknh������2�4��̭ߟ!Il�z��D"�(YK�pp�3C����s&�^�G�3"q�:y�}��gGUY�t��+�6�����d|ƚ��ɶ�7�' �Z�ե ��X��M��������X�;��~����f~���UO���K���rGr���Ø�������Й=�T����
��ƧڂΥ�w-�V������]���<����x�K�ؙf�C,u��Yt���J��vژs����
%��'�&�'r������ �\A���H�O��ܟ���y�VZ�H���'s��eb~�҄(�i2Ք	�]/�〔��N��J��	+���F����n��a��GB�S(ڤN�+=g��\=\=�,>2�I$ؘ�r?�<���կ�[��7
ZT�_�0.\��Մ�QK�;����^���e�'T���4]w<���R�I��*�2���B�YWIVV6�]�=.
Q\�Tⲷ��������]8������������k<���<g2���^h���S�s�?�&�Q�X�BTal�V_�@�/��B��7�Bm�V5T��V����j�x\�0���~�W�kBr�;)NL\�.�8 ����(��_�r�R̙�|3�rQf�P�l�������Q��;s��M��m��@��S0]}�F�y�d�W!|p7���[fK�&��Hk�NW�8֩���q��F���?�~G��^l4�V2
���gĳ~cx�"�,-UVl��_o�	J�xy�����x�M����ۢ[a\�r@�����j���K����1	�WQ(�Ux�rD�9 =��#Fn�AT�����3�U�M�3�6��C38,-|�}�C
/k�G��)f/�\����V1�ic���3k���Z�on�؄��E��sw��B���9SBpQ������B'Ƨ�z����wqR�1����E�m��F��sZu�+
�C��e�&�{����@�%�*�v�2�7Q�ۓ-ם�x�G�kFÁ��u��N���n�����w�t���3�ج�����M
����v~7����h�Dt�����R��m�T��^a���&3�%*܎�X�Y�T�
��p��+.MӀ�b}�%�צ���� %�8Hq��-M0���ׯ���U� ����b9�}������Q�w���K"$W����3=8jԂo$�S��=z�����D���5���vҺ庙J��T�̜g��뺒	S*�	3ޤ �ѾP�~.Ge�l����a���h\��)v�%��ѾO��/@l_�{L[РU$Ǐ&^��`ԩ���'��e�� �z���	�恗��dC�����U����{{o�ʏ��Z��������e�M�`�&Ôw�b��#DY	�[Ԏzc= ���A�Ca��eU�H� (EVV��[϶���]s��K*MQ��2m�������� p��l�t�)Cd}�ĳ��9$\�?P�\� ϡ��$�0$���WMxc2��B�G�ݗ�Voqm�`��)9�>׭ɒa��гY��R�E���@lT�Q��Sᜣ.)�����V�6�����Z(�ic�1/�}� S�,~t2Z�dL> �;�}u�6�)�^S�z:��Uf^f�V~c��.���
�_��TW~�<�ő��4D���t�F�r���ǀ���on V=�R��=������@w����4};߆���h'd�"`����uk��D^�_��F��n
LJT~��
�W�aO)��}�I{A�4mYn�4�kSKH�G��T$��!4��<���݁�c+{�����֍Ko�UEn.O�Y�p�r�oeNн��m|�:(I��Ss����~N���Hl�!U"�!�V_6��/Y� f7���x�x���m'��"��P���Y�y�JX���m�����o�}!j���0�U�ϝe#ǽ�	�F��,�+}�7�@%�UJ����_���1����%�_��,1�}9$ӣ�W^�W$��0����FNV����yOi�O
�=­6��7O�����#N�d���K��-�N�i� ���n�,>RT�U]�p,���R���Ud>w�o�!�:�Sh��5�2��s��N�n೜"َ�Y����}�CB$l��7�',h�d�.�z7�:���m=�r���/�;�����] 4f���V
�:��5��o��yg�n�C~���)-���_�P|V1�M�#4�b�|���)�q :%;WQmkc�j�׼��*Ҩ�8�c��en~�/a� �-p�o�W����>����,�6RU�i�㢋�
3(���Z�<
;Q.�P*K$�TDZH�-��X��u�$��;�IC��Cȧ�+�>Q�e��x� T��bu�C�W��I�p�6� �wl\��7�5�~;�(o.�*��h$�8��[�Z<��}��[�jF��`����H���S�b2��6e�ͥ���;�!O¼]���%o�Ct��;�a�#�C�.�ӕW��R�Mcz;�>|�����v�*�`g���{�0B9�+��i/���U#m!
��T]�i^�_a��-��[S�󃱫5e���2D�)#E�x��C�̇ٙ?�_΀E���B"��wqf]�@�a� 䑾!��R��¶d���K.�/1R�n	untka��י�N��,#<d�D��8�(�(�u�#^o8 �y��\ʈp}���K����Ɇ�����ci��w����gE�8���ϫmw&��]�u{�/\����;�S��'�.��l6ni^	"�_��Z_�j#��f�v��a��@|׆�w6���W6�c(��`cł��~\s�aRY����͟,5���O9��Zȩ��6p�P4�-�.l�������)T��T��l����S�&n41i��6�����" B)������DL +l[Z.�(Q�9�3�Ҧ���+m�>���� �k�%��	���~�`�F��S?}&�{��*�W a6�Y���"pU���f<\�M����it���@��,�ހ�ctkN�s/�(��H�����x4�PE��r[��V)M���kT�5�ڳ�w�[����&*o��v�z�	;,��G���'X.����@���8��ݗMoiLD��%�ڴʞ��~$[Qg�BN�3��[��`��`@a��D*�l:�g<S90N�11B�����:l��m���j�3�"����Ea<��������+E���o�m�z��Ŵ���c�b"�5��!�ϔ�C#�2�G�8��m��4�������Ո=C1J�l����,<�k���g��G�5������B��0r ^mcH�4匚�^K��wi�.r�ȏ��|�y�qJQ�f�O9�������m�B�S.?��20�xhX�5��h�JIP�RɸZ��>������,ߴS��ڈ��%��ū1��2{�� [�}�o�hQؖ��ï8w��� PpG���y�,�S����kR��/��� #K�^��0e��_TN��5I�~�*ѯ��Oo)�\��-�$��V(Y���A>��L�-�(�hN@\�b�'�_�g+�G5$��}�!���T��Q��aAΦ˳��O��P���"';��$�6�;�"���WIg2�B�5���:�|R~��U�6Ҿ5�@�B= �(��9 9TP���zO���}>~n�bD۳b�����3�	�XJ�m~���Bu�������܏���S� 7я?~ ��D��}Z��iݨ�7]�_luZ7^��bYSB	�q�}ħ̼��!�H���68L,P.�{�$F*����lq1�apQN���\y���W�����{<��ޒM4�Gop��v���V@΢̆��=��{�K��^�U��	�h�%q1�3@�D0禡��u�PE���i�s]b��5_�@�{q�&��d�':���3�F�7wT,R q�s�>�r�SE_��^f.�����C�
*y�{�����e�J���B-�l�j����U���^��:Mx�x���@�q`�p���p	��ب�f��T��9.�����@��'+~�S�ɸ����`en�K�Y�c�R�o}���2ے�֞o���c�#��;� g� �=!TޜƜr���Q�����O+E�Nc+����������y{�̀b~ǥ�i⧗����O]~� �I'�浫#}�K��pG���,�R���T8��u�c
核��d�7�0&�&#h>T�WJ�QVÕHQ�k���o:�o�f9���p�=
ucqW�z��.d~՜޲���!yI
j�W�̞v}\֑4(j��{�{ ��}0������JR��}������m�Pż#/�%����a�h�#�8h�f���~q��Y�i��B�ו�*�qjD�����5��?������h�|,st{�o�g�予�gi��iq �
^@��g�6��/�I�Ԟ��($���l�rDB����wk��"zB`e��kT6"C�b_v�+�ji��x��W��ރ��	҅Sq�����m>N0�B�¹�!E�o��ϰ�����ѦO���hG����oÍ��HB^�e ���ަ�*O��y��;+Ֆ����\�oBXQ�&l���o��u[X]�j���կK�l����՟�$�~����n8 	_�,�fY�%�i�ܠ�[�`r!G�������b��W�)�"}���M�GS^�� m	O��ڡY��Z�Gc;j6�������z�]�[ Ӛ~��HIH��3@�+du��Z��s��2��N���gs�l�9-0�D[ b �Sع�J2��z�i�&2Ö�7�}�/8z}j<�!�^�Zl&�
x&�bU`+j5��J��^A(�����P��&�<6Y?�)fc�"Z7��$��H*�%��u�M�,h��;�B�����O��w^M��:cm-}�NFY? .ŗ��!��2��D΂7x���!��>lb�fg�E�M�aN��j> �n1p�O�b.��njL�b�����Ή���`ID��^ ����6�nk|z���?���~�� ���jY��i���|��(2�a�L�n֌m����5��oL+'?��S�2�~.?�|�.c۱ӱ�Z��;�B��z�:�x���iI�h�Hv��]S�i<�3����n��J�g�_۾<˾�V&p�uϐZ��&��C'����QO�)�*v2�*
4*W����m_�GK���'�mD��	��!p�� ��o��DM��,׷�0g���{�;���5��z�r\�(�����m�>� t1�H�1�#���II]�a�̿�-���Jo
B/�O����I;�)� ���q"����M��&%8;ຬ�����{Ʋ�ݑc�᧼{/���i�\�H*���Is����6hD���fI�>���tK��G���@��&5*8�����Tl��	�5����OR���qܡb�X�|$?܄�ch�:&b@��O(��P���BSWAG�0}�=`}�7�I���p]�ӗ` M[���Ƚ�w��<�����BGJ�c� DYC.�9d�'��Agi��dy�~����:��5�'�$ N/��-n�C��S������ӿ�U:_�km�����Ƭϋb2\���Pc�e^^=�����8s޸ᒾ=�$�6K����.���2䝂�k*ǏE�ԕ�����>��i.�]�`@�;��r-�籱���P�a����P%���鈦�����ݷ�lx}�������`���M<t��������2��5�4���M��m�䓭�)(���~�j�4����8�z.��,D�l0����~���u��5A9���{��租ov�Ɋ`�[jlL*�^m�^�u�S��×|��}��ڎj.�[4|��剆3t5�/g5JЈ=~��)w�� �W�2���^�a� =8�\~飾Z�6�_���j~����n���jIF�^ntu�$�>�a��=�9c,T$�I1t����ChOĹuӂ'�p�P�[� $.7vl^�Г�f�@�	�7@U������r&��]x�^ّ��׊ ��g�[T�ޑ�!_�W�G^o�<�$��|��۟�j0�����Y�?r^�ȓNs�?��m2��� �T�k�@pB5u݂��Pcx�l�ӂ˭���;9����jTʏ�T�+�i?n,?�ؘn��D�����W�mia:b�k@G��k�C�:�I$b�ԃ��/�p��x�{�/�$N�*��!�S�F�=l�a�,u�mӲqiCH�@�6,���ƉXI�~�O]c݂}�P��2�`��@%����'�,�NO�����B瞚	�W,��;�cA��e;�*��(?��^{�t�,�����
��Z���|��}�iʱ�����מ��]�?�X�X�wz������V�ۡS,.��!XdYǍ*пc��}�A,�$��������a��d	�\���[��{j��Z�k�O�9$5Il	�A��D(�'���O���������3�k"E���>�l?1��4�x�0�<�Ŵba�{��e5	�ϗ�GE#�JC�_��[��ׯ�U���=N���~�����s��`HN�خ����,�kp�ZȜ����W���cC,��&ǃ��V��g�E�39�2eZ�)9��{	���U?2��s�N�j���M��	�/�=}� �����vʹ��E���&0'�Cg>��D[� >0?��{�������u���E����)j���o�k̄K ��Ǳ'[������,���} ����&A���5*��4Zp�i�7�0�y����K7�/v}ĝY�綗0�0�T�p#���P�n��}�Ņ�����(�N6��| 
T�����/A�*\'u%.��~ֿ��燍��0E.�F��mO���ҽm�~KznO|�#��K��P�H�V|��o;q>p��c���pkpR��[�Ԧ�(rEV!�.��V�ɲ�bq��[�CkPC������ؑ>K�|���_�QSn#</��q6�"~�;7x,�;~�x�C(�`�3�s=c��ƪ�8ng��w��!իx9N��	 �D����夒�-�1�ǹ9��dam[�F�f��L1��`	\�Ҋ�2���Q1f���A ��Z���tq*��K���0�B��Հ�}l4�<�u�ֶ�Mw��ϱH�=��M�P��C�}<^��@�2��C�:����P���_�}X<�8�[�ECD���Cp�o���íӚ���^o6Q�6��UHU&
녞yC4)$A�͇��-�4�gjSO5/Mn$��I���<B��|E�h%�\;��jA�����8�bT�yu�0�I�*��:3���Ix���8w�c����7�۾����kP��Vz�3���d[���]z�}��|�B��}��������%���%U�H�
��ܢ}���V#A�H/����Ku~2�1����؎6���6Ǹ�DY�|�`��ߕ�~�Gt+�\��'��M�����<�eq�>��!RMg�_�&��ά�h�g,�M+����[{�j���90����$����|J�M_ aX8���s/��	��;/K�R�!j�˅[~�g�0��̝�b���7���{T�鴠R ����$sf��~gu�w_�}n�wQ�{_�'U������tciB���5ĻR��,)����iߕl�Oݤ�f5�k��M�٨Z8l�\��X��s���o?�j;e�>����}�ͦ�Ô���,6��H������G1�rǲ���c���y/[ih��,��N�\����� ��#v�u�y�}K�7�7,��U�B
1���v��è�+j �gZ�dȞ�y$3�lz`�,/�k�[	BP��^���L6z�`��7�Kw�_b+�CsL)p&2�Q�i~�z����l� p���G�*�Ɣ�L��3b192��j[M�9�aou���9D����\�߇�"��7���4����a�y�p�Z�������5���~�,�VY�Xpg�c`�˖�1�Dy�g{����-/.Ȱ+��K�dS-��/9�Ӽ��̧z;��ΐv���-�I�7qӮ5ۆ�������w{�Т<	Yx�8���,�Q����/���&=���Nж���Zy��wt��Ck����7t��&qXM�b�,�lE'��vTD�{?��Q,��h`�=�.	2��*L��S,�}i�|3��}�RY�U��|�Dm���*�)�o��	4p�}�J�>�yn�L�E{��[�l������
Q{v����xF4}6���Jƞ"����#%4x"����37
�=�U����뒏(2FJ1TUR���[�wf~�j1��,� F,���N�
d�`��/�5�߰Fi��>�3Aݣ;���G�RZ�����TxA��	�������VQ��Љ]������.C��_�,�R;��E��]�8��׿�ݘ%���v׻�`W���sG���2C���)-4c������}s��5���t�Q�n�a��vN��^�P������u{��/���l��8�N{P�-��d�Z�yc6����^u�@QY,Qw]�l,���d�JoC����aϐ��Yx���@��`iYCXWl���9�ע;N��ʌ�o�ORƷ,F��/��%�"U�=4�bz_��C/�<:��<o�f�k�E��S;�y�)�ϣ�3�B".���,��In�6�֓���L7��忧�Z�!U"撺)��3;�5��I�c���c}��?w1+���&�ɷ�8@����|�0��',�+s*9�|��G	1V`���<b�	�D%��}G�)ֿ�|��I���B���ޮ��|������C؝ k(^�s�������c��H���tĈ�$U ��V<v�dhn���+�w0-��S�q��-���K�g6ש����J�S�EKS�����L&�P��mL(���^/;�|l��`�u�h��]¶_a�!Я��{E��{e7)�2�H.��{/8��q�'����z?q��~ ���+^�[��c���p�{�,nV�b�\�|�R@��{2�E�V��X�V�z�W�Ig����'?3�Z��\�h�˷8rC���Mnz\���c��$)����:���u��rv�9�F��(��=�C��b�~��Tu=k��7G���&Y^lW2 �V���'h�6	8��A��#������N�K�7���Z�I�<ڔ������ T��o������yI�#K[�Ҳ�~a�6щdQ8�W�B�Tr�:NQ1�sC�X����������H�6.����"/�:�����j>&�=	~=�'W*�_�E�W�z �Pʧ�|7��VUt��T�� ��˙Zbp�%R����Ӻ�;��-����sJ��:�:��4^T�6Ꮜt n1]	7��M��: �����V����%�%�:��������=Xe��J���*bH,��D�p]J�K��Ñ��P��8�?�~��OԒع�����I8�ӈ�zo��� 
_B-�/7Z_�kEF#�����B�v� �jp r�HIj�<T5��؁;�7|���{�dhc^�@��,��薀�g@+>�QI.|��n%��9"�)�$��c=d42��z��(��1�
0��7�	���7;m
�?/C�|:^Qj���&3F���$Y��#�ǡz�{�ξ��J�Ӽ�;�x\��X�eP�\�"��#�pU�6f�,\��: }�Xc'�S������N)�Û�����0>������R]�룥T���{ۓ.���_K�r�T[6����BR��Sׁ�̢��X���W�	#K�r�>V�����^{Ѥ/�atiYʛ'�ܿt��/�������>��gd�i������Tp��8��+v 2�����&'��+�>9��ڸ
�8,!MI�Wf8�>j��Szwњu{�N_��ɗ��{��y#s�iz�GG��+-W~0�"i��Q���8��N���"��@G������n�o).Vx\U��%�����F�b~G
����j�v[��:̾˱��_9�o��)�WH&���P��|���0](�C�|0���>ܢK]"r�/sl��g�m�⇸a���H�8UI�
��@��<�u z2Wb��G��CsE(�c������?V�i��y�TXbظ�.��?���:�5�b���sJ�3$��o�>�I�3Ht�?��V^����}�6�S�����C��ŕJ�^&�P /gY�T����b��Y��<�a��m���U2l@xc���pfNP��c�T*��Ϻ>J�f�/�h�t� +Lg�H��|g�B���^�e0_��G^���� �T3�K�,��x��HJH�4;��V6��M��~Y�3�/�`�S�ZB�`�귵����#G��0�I���A�	\�p�xh��$V�5��Z�rW����ǿ�3��߂YZ�U.$Hb�y�����nU8|df��I�N[�l��(�Q\|(s���Nr��j�Cˣ�������n"���T��P���z���/Vԕ��H�/�
{�����i�!'B�e�H=�lJ���)ǌK�t(��}�2�j�:�+�tW~��~��`�����BV+)`rE���S��&p��R�1BŶf�;hŜ�13�{tI��2��7���1��ؕ�
c��Po����PQS���}���=���4-6W�`q�07d�bX��LB9�W�tޒ-2�WW��)$���Bh?:aO�0���xyy�)l�S�[��e�y�!N [�b=`St��ע̻�GvV��O<��X�	Y0[pziR��0S!�b�Gq��M�H"���4n���$�h���C��lɕpN �jR���Ү��(�?fʃ:��oم�0��ョsޗ�&'?೺t�/�=����e1���~��1g���_&�$���͎̒=ٲ��Xk}Yjtj�[.�	)g~�1y�qa��^÷ Q������i8p :ӤC�<u-���y�z ��tg]oz2���9��Ԣ�H���d6j�F� ���	�����3������c�x�e�*�|��TT�k����p��Υ�ꄥ��,�W�4�+���ĐVfO�yq��;�Q]M�|��E�����:"L?�=��[�`+�8�\y
����*�[������Ǽ2��?��(�`�~}��n�x~����i�ԭ>W?h�˺s�>O�5%�� $� &%���y#��IqGy5��Y��a8��~n��rα���y��2�Ov Rh���	ce7N�BE�i4 { b�s(7(�)�E|�@l�>\�����?���v	��{t��	�6,��b	�Ş�	� �J�P���|_e�K��*��iᯍ��_`�ߤC��JfO��H
���'�<�n��y%
.q��0cX*��v0~�W�9����'u�>�^�����g�gq���j'�]��K5Ԡ�ӎ��m�/n��س�s��S�,.3*�?꺸7[�����(�waEY�{��;f���0�!���C9 ����Ȫn��R��w�-��}3a���C����6���@2u���I°���Ԝ7�����oa��f�{&8��O@� �g~dI��Y�3�e��s��OO���j��v�c��9Ö��o�\�? ��:t喞h�����.��v9�}��g7���������������CV�M|9�!�E{FUn�%��u��dt*�������{i��n,5I����Kl�k�����=è��V�Р=y����p��?����J����F@�����-x��E�f3ݷ-Z�qP�s!"+���]P/�~���k[[�s��.�cS��t�K��w�B��*�< y{��d������
���W<|u�(h���ч=�:��U�^|�p˿�k�T�$�|V�J/Y"��.U0�PI�'�v�P���	U�j�t��Unz�!G}"��9 ��o,�J;�ɂХm�[�XOn���I��x-�� \>yԽ\]��?���O�v�hƈs���`fj�������!@���Ưb���s��bݖ�E���_�Eh)f��в��!S,	�w?���5¾�@�!��&~A�: q�i@$�'4�d��t,�_�ZR����)�߸Nl����bN���i�X��t�����V���s�&ǥ�͈`~��r�.hYˎI_W�~������oh ��0�l(:�/N��S��2&��cc�C?�ߪ�V:сYRf�6�ZY�ksy�@�u�=B�-'fm���
�����r������6~��2L)���p��+�}�+��)�~��Aw�'O�jm�h��� �/�8k� TmE�Br�dޫ���v�}�fZݽ}�z�bϑFӻP�XU�!6+6�=�l;�Ģ3�gK�mV����u�"�����c	�z`g O�3�Ī(��Q�V��_��c/}:�9�g)��N����<�������u�Zۮ}�^��X$����&��5F"x�1&�P�&���'w�����l
T.�
߮��޴�'I�w�����K�3l�C�BߘS�0�>���Ր���^zٟ���NWtu�'3���V��T�^1���xB<r�c�i����0�
_g�v\a ���I����VAdE���	��Of��Xt��;I��J�ʟ;���.I�{x���-�{�=����虊���]�0�)��j�U�GZ�L��s���&���������;aDp�vc(�.?�Xɠ��+���z!JR��r�%؂{8�}Mb�i�fn,���L��lF0����l��O��q0�2�lMQ�Ҳ�}� ����-��G��T��$�t�e��]�W�������<B�5l5)���P�zCӾ�<��9R\�!�N&��O�������s�25U�*��j�����,�B��8p�!����b=2r�G��ђu4L/�K$/Á�a	۾��%Ï9�6O�}R��:��J��2|���O���`���QG��6g9�;�5��/��r=����f��<�u�K�U7LC=����ƭ����,=���0O�K��K�]�/w^���+��{��� �,�qHY����.u�����*�-��A�2���t��⢤�#ժ��l>�L:�P��n8x��!�O!]G>ܥ2��5$�m*��A:����Ց$� �W��~���P�Ю���I��x��х���|/g���Dc��L�D->� �X��'���8��4{��a���_�e�&�vJx�������y�׀��`��˟ 	p������4J����L�![�5�Iُ�x6���q�v��{���3����f~���A����s�"~'"с�9[~ɽ0у<XŔg�k��+|~��:��QU�5�� �o7�K>���>�nf3���,�Lh�����������SW�wY�I(W�5��@�*PL�U1�^��L�QSw,�9�$�5���ď �|��G�Y'#*����Iy��;9�C��L�M�mR�֤��N�^��i�H�{]ej�h#2L�	p�O�"�5�H2���2W� 5��[��A���+�0,�ݙ�������S=����1��<j�O-&���		t�	S�� ���uX}tߴaHN��i��]X����Ҹ��V8YF��݉m��m�.T�o�H�H��k��D�t�Y��Z���Q�����H���~��,&�.A���ij�Z���z�C0v҅1�m�ek���˂�#�dp���7�vb�8�r�׍�T����0�!o.꭫6�%v-`�0���8�jCV����W�Oѯ%����i����(����Ռ����
��;2|�~��]: ū* �Q~Տlh�����V$;�O�
Y�O8)Ĺ���4>h|)��썌U�-���{_'9YJH�>�����m^I���o�a���W��Mu0jE�fGŴ^'��[�$�pTA�R]�v��>.\�\��gq�/�b��6�SOP�������њ���8V���	�I-���Q:���$s�ױ�`h^���6�d|F������i^�T���q�� D����2������i�V�w����� o���R�s�I��rEG�S8q��K�φ�vx&���-�NZ�M�C؟���l.tSx�`��<�ʰ�o_��v�I�9&�S~g����o��~�}�s��*�!|�F=�O�URhҰ�$����a����U�V��,\o���;�,ffR=6�5��z
�&��..�t�d�
ʕ
�H��b�.¸aԏ����9�L%D�g��h��Od>k`�׎���%���Q�tG������X�����/����`=�
��5�.unF�\�lױw_��	��?p)@�g�'�N��k*G�l���g���?Я��m���,� �@� C��t���U/���`q�����B�7ͼş>ұ}���wks֌4��ڦ�d��=5�к}2���'ۡ�w�/8�V��ji6���5�����'�2&�tKpi�_"\�$p���/�Cw b[�����`���P�u�mS�Oe&����O�<��N���V@��F�q�k¦�tQ~�{�	+�&�� �X������:���ʙaW��PHE�=���V��5v�z˭��}�V �˕ǌ�;}�g^��ͳ�JR]�n�nc�T�0.�Yl�u�����"�V4���^�s��,:��ph�$ɳ��
�;&ZQB���y-�u�A�'،�D[�t��a�.͜�}_KNݐ����b�X.7e����=Z�ۋ�Z1�+�� ���7(������Փ����q'h\��$���3���$?����;��L���b%�Ź�a�w�˯�����Q���v[p�7�86��IUz�1�뮨i�t$��\�RD��I�u�PN{��n(�2d@�I��iM��X��:�[��P�G��x�1"?�4ź$����ט�(=@����Vt�����������3f�r�a�M��kVǡ��w��N�M�-�J�
�d�]��P8�5 Fz��(��{�B�ɚ���֭/g��S�;R���).m�ɻ�a�2-<6s�<_�����_D7�ҭ�|��I�Ȫ�(���9�����9��M���DsVZ�M��g��?X-΢u�(,;��ϟV��I��ÖZ�o�;��|�.�d��wL>4�u tJs�����sr�=�{�X�e�$~���j/�I��cj���w��{�_8��%~,޸�8�g�]�WX����!��T9����Ҹ<������]����:��9��K�8�!ԍv������	!�C�{�5��F���v9[�:���S���U���I:uu����-ID3Z�	җt�碿������gA2�3�LpGڍq%*�B�����X�N��H��èj�P]6¡ B�o�)`���A�2�)k˄/�����w&ޘ�"k[���C�-$�r1mw�;�$s{C���|�?��/��#5���nK���u�1�o��Co���"[J��F9^ْ���S�9�s�q�)i̐1>�y�B�)���w^8s�F��7�\����V.�=�B>�g�uΦ`n7����9�s;^���?􍉒�|�K�j����]���ؖ�À�����<#-8?���ɍQ0O����{���o
��gگ����Ń��E�@.:_I���\':�p`�O��ء�r���TՍy�������p��Ϣ��Y܏7;-`g�j�HOlt���f,/�캘Tԙ��©9G�j�
.7ҍ�V>�l�N�
AK��i� �Xb�Ի��dGx���G����x<�Uݘ��OJJ����Xw��s��ǅ{���ҟn�yE�3�!}U7�<��L�Bq��T`��]m���UMM�j����e{^:t^��ˍ�q����Z�L�%{o��)1�Jk���z'��ۤ�xL=Y���ɒm���8ʟLV/�!����>7'�9����u��QZ��bi ���A�K�S�XpG�x�� )��1�m���LuNe�G�FэB�2'I�ʿ�u"ܶ]�����3�_ ]෻&�x��i;�smu��뽯���=^q�oQ�}��3�=��
�-�~�K3U�[���(���f h�ɾ�4ث�<f�W�JcD2�6AY��n.^s�����T���1�]�[S�7�-�kcU����y�n+Ձ'��bl�<%�sf��:��:��	ʏ��;+@��|_J���.���uȫ:����b���Wqԋ\�y% c��n��,�٪��D��i|���������Փ**'A�ۇ\͐g� T�K�f��A�����`�gs?qh���Y5?����q����T�(�h϶uR��g#�f�^��}�S˓�E����}b�q�3V�0n,1W��כ3�%Ov��9ߦ����} �f�L���Ѓ��jb 򨾩����Jvxɩ��ή�L�!\�����"A7���y���)�U�����K�!��s�'RO��;�}.����ayH��>�P��o.��Fx�Lɘ��ƥfP�d��.=}wk[˶>� �������>~p�L�#!�]wK�2'�p��zI�^�j�����,��i�Y�&���=��)�WEWa�xA���5� ߽�g������Y�������~�W��N����X2�r ��g��MC]<Q_o���s>L_���w��7]r��RI��^Z!� 󘒙h�^ٙ[zCJ}p���ڋ�LR����u��wV4�p�H��1ň���x"�\�C�_�l}�Mqb�xC� e�nN����o �
�vn�W�~+� *l4��W��e3?Y�����ɇ"t/W��X��
�@j��/1���%tVD*d����Wݻ9n��Q�'Rd�b��s�VN���'1���W� �¿J��ź�@I<�ݣ2_9Lt6�좽�|!x�>*��Ǘ���8W��ʤ4{j�/ڃľ���~hz;,���Z����ht�CdnGem�)�f����e�	$c�_�w�� �~"��>�����_�$�߉l�.��U��6b)u����idfDbrr�����Lf���
6�~e�T�s�'޿����?G�2H��Q�����/��\f;�
j:�?w�� �����K^�Ɖ�^�5��\�(��6�R?5�%'�	��_��RL�B2�v��)���_������?m_��Xu�|%����0�.����	5�df��H̻C,�؈� ����Q�r*�
r�j���c�5#Y�={�����>°��MH�T�jbu���A�'�_�'�G�k>��5	�sYA�xH�����y/��G�@��5��� ��� �n���py��|��B�YH4�x$#`��������-��� �=��v�|q����|I���`�if�Xm�� vm�a�c?��xEW,���W��4y,��gX�_��:V�{����������Ѵe��1o�YQb
��!�p+�����O�'���@�D:��9�.,�V��Sq��t#��O���;���'�6����1��F8��DY���*Izʄ� � ��}{�_�O���O�����)<���k;�O�B�����I�qM�h�&F�+�87��,���VRr����ߜ���j�k�k|�~� �^���嶳�3K�T�\^=�潅�i%]�X���ҿVj�#��W��!�K;��b�IH��Ǔ�ֿ<��Z� �m�i��>6��}?��Mrm>+sz�Os�Ѥ�<,Й:���v�v�^��?�������k�~4<�w!c��(�d�w��1���y5��>
T��OF���w���������K�j�,|��w�ӼG�0k�#Q�4>+�1v�bcx�2GA�⿧}+�� ��K���]�.f!���Ic����������N]c�j��>���ZN��\�qޟ�$�D �.;�8� �{ѿg� ����K��.�,f%����t�p׆L`��~4�CW��[	U|*>�� 8O2���(:z?5�����ľ���1xx���u��
4��������M��YxW����n��ii���_�W��b��U�Y��J/�˨�Fm����$�bY�iN�}�*�-~3�i-��@��S�v�����l�
���//�dy2���v���?㼿2��9��Fϥ��?ً�
��m~ʚL>����hO�l�71)�^�aG��^����}� ���ɼ#s�X�~�T�?�]��ҺGvߟ�N�A���j�K&r���?�U{G���g��a��jK�������s�B�f���dr�����8��G�e�y�յ�Nm[Rk�����o�I�L�.��s�`��A�&����b��~6i�i�_ە�������bI�~�C��q_H�>� �����贏�>�_��.��S�$��l.ݖ�)�?7 g W���f�̩
.�1�
��a�t�9�5���8h�xc�,�����'�3��PK   ��W����  2     jsons/user_defined.json�Xю�6���_#��\����4���k�
ɢS���v� ����%�l�q�hI��V3�C��>l��r�����&.�.6�b�O��Zire���G����?~��z7���}ۭ/n��.v��⅗�j߮��`���_��ES��F�a4�	K�BU�[jt	�[~���;���r��㗽��vѷ���F��x�.2�զ{+�6m��[�g�g��ݼ�nVՇ��j;��2��Ђ�{����X��`;��ڿ����es��[������W�J� i�B�!,�5@$ϴ۫n�纗՟�tU�qX�����qxL�@1j��j�5��3�� 8)@u����~z=?�O	>� =�ɒ������ <$�ޢbg�.|P`]S���������^޷���^.��M�w�2j/�݉6���~x�#��QMk�K�)J���*.�eU�YR���^�!��y07�!����Oאe�<�҂����:��$O��{��9��H��VΑ9��F���J�����`y6CR��\_�6���5؊˪�TR��ƹ����#T�������6S4��@֏��<x:ύ���@h�X9$V�-͏�0e�!e{S�Xa��	S�|@\ :��I����x�\�.M͹#s4C`P�
����Tw^A	ؑF���(��8��ǃ�n�����u�N��H��sP���� P";Y �4��A+����1Ny��nP�l9%LB��?2DƦ�%ą�%�%�M%��g��S�:�
��A�A����L�S]>� S����@��s��z��%:�%���ꦌ��&�8g�||F���~��H�!~�	'����̐e�$6�ѷZ�\@;|HJr,v�㏘��i�Y�����,�t@�`�#g��� �2����~DA�ǋx�p$�w��g����#�,�+'f��"O�g6�S}ޮWUqSuR=��!���!�KZںu��W� j\C�h4>��.�����H��g>]�"!��`,�	Z���0��;�?���#{n�G�/@���^�PE{�M�Q������J^�$���������R%>��IN!�vNʡ'w:QXR�Di_��d�r�*βs�Y/&�aN�ϲ��-�`x�+�
��9z+������������H)>��x�U�xq�T�]�s�c�A.f]���z_:�n��Ϡz|�%�:4�n��w����Ca�, ����qD@9��T� J�M���1���o�?PK   ��Wx�D��,  ��            ��    cirkitFile.jsonPK   ��Wtk��  ��  /           ���,  images/0732da8e-2e31-48ba-8c11-1e28d7829515.pngPK   ��W��S(^w  �y  /           ����  images/2e36d9e2-369a-4515-94d0-1575017f862e.pngPK   ��W��Ƀk Jn /           ��b6 images/8d0bbfdb-2662-4be1-b50d-e5d8de487479.pngPK   ��W��(��� _� /           ��2� images/b4c55bd8-374e-45a4-aecf-ab43f4af1abc.pngPK   ��W�6U�o � /           ��Bh images/b829761f-344b-4f5b-9b94-abe91c4d6d49.pngPK   ��W�iҶ� t� /           ���y images/eea2c8d7-d880-4d78-8cc7-667d8a2c86d8.pngPK   ��W��s�2�  |�  /           ��B images/fb2015a8-ad74-4a61-8d66-2e77d7201afb.jpgPK   ��W����  2             ���
 jsons/user_defined.jsonPK    	 	   �   